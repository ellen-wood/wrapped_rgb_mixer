magic
tech sky130B
magscale 1 2
timestamp 1670930158
<< viali >>
rect 7849 39389 7883 39423
rect 16129 39389 16163 39423
rect 17049 39389 17083 39423
rect 17693 39389 17727 39423
rect 19533 39389 19567 39423
rect 20361 39389 20395 39423
rect 21005 39389 21039 39423
rect 22477 39389 22511 39423
rect 17141 39253 17175 39287
rect 19625 39253 19659 39287
rect 17141 38981 17175 39015
rect 24225 38981 24259 39015
rect 7849 38913 7883 38947
rect 16129 38913 16163 38947
rect 16957 38913 16991 38947
rect 21097 38913 21131 38947
rect 22385 38913 22419 38947
rect 8033 38845 8067 38879
rect 8401 38845 8435 38879
rect 17417 38845 17451 38879
rect 19349 38845 19383 38879
rect 20913 38845 20947 38879
rect 22569 38845 22603 38879
rect 4997 38709 5031 38743
rect 16037 38709 16071 38743
rect 28549 38709 28583 38743
rect 8033 38505 8067 38539
rect 22385 38505 22419 38539
rect 4905 38369 4939 38403
rect 5549 38369 5583 38403
rect 16405 38369 16439 38403
rect 16589 38369 16623 38403
rect 16865 38369 16899 38403
rect 19901 38369 19935 38403
rect 21281 38369 21315 38403
rect 7941 38301 7975 38335
rect 22293 38301 22327 38335
rect 28549 38301 28583 38335
rect 32781 38301 32815 38335
rect 5089 38233 5123 38267
rect 21097 38233 21131 38267
rect 28641 38165 28675 38199
rect 5549 37961 5583 37995
rect 19809 37961 19843 37995
rect 28641 37893 28675 37927
rect 34161 37893 34195 37927
rect 5641 37825 5675 37859
rect 19901 37825 19935 37859
rect 28457 37825 28491 37859
rect 32321 37825 32355 37859
rect 29009 37757 29043 37791
rect 32505 37757 32539 37791
rect 7297 37621 7331 37655
rect 22109 37621 22143 37655
rect 32505 37417 32539 37451
rect 22661 37281 22695 37315
rect 6561 37213 6595 37247
rect 8401 37213 8435 37247
rect 18521 37213 18555 37247
rect 22017 37213 22051 37247
rect 32413 37213 32447 37247
rect 8217 37145 8251 37179
rect 22201 37145 22235 37179
rect 7389 36873 7423 36907
rect 22201 36873 22235 36907
rect 20269 36805 20303 36839
rect 7481 36737 7515 36771
rect 17785 36737 17819 36771
rect 18429 36737 18463 36771
rect 22109 36737 22143 36771
rect 17877 36669 17911 36703
rect 18613 36669 18647 36703
rect 17325 36533 17359 36567
rect 17509 36125 17543 36159
rect 27905 36125 27939 36159
rect 1869 36057 1903 36091
rect 1961 35989 1995 36023
rect 17601 35989 17635 36023
rect 17693 35717 17727 35751
rect 29745 35717 29779 35751
rect 17509 35649 17543 35683
rect 27905 35649 27939 35683
rect 19257 35581 19291 35615
rect 28089 35581 28123 35615
rect 27905 35241 27939 35275
rect 27813 35037 27847 35071
rect 9965 34357 9999 34391
rect 9873 34017 9907 34051
rect 10333 34017 10367 34051
rect 27629 33949 27663 33983
rect 10057 33881 10091 33915
rect 10241 33609 10275 33643
rect 10333 33473 10367 33507
rect 27629 33473 27663 33507
rect 27813 33405 27847 33439
rect 29469 33405 29503 33439
rect 32137 33269 32171 33303
rect 27629 33065 27663 33099
rect 31861 32929 31895 32963
rect 18337 32861 18371 32895
rect 27537 32861 27571 32895
rect 31217 32861 31251 32895
rect 31309 32793 31343 32827
rect 32045 32793 32079 32827
rect 33701 32793 33735 32827
rect 20085 32453 20119 32487
rect 18245 32385 18279 32419
rect 18429 32317 18463 32351
rect 31585 32317 31619 32351
rect 32137 32317 32171 32351
rect 32321 32317 32355 32351
rect 32597 32317 32631 32351
rect 17969 31977 18003 32011
rect 31677 31977 31711 32011
rect 20729 31841 20763 31875
rect 17877 31773 17911 31807
rect 19625 31773 19659 31807
rect 20085 31773 20119 31807
rect 26433 31773 26467 31807
rect 31585 31773 31619 31807
rect 20269 31705 20303 31739
rect 20269 31433 20303 31467
rect 20177 31297 20211 31331
rect 26157 31297 26191 31331
rect 26985 31297 27019 31331
rect 10977 31229 11011 31263
rect 11529 31229 11563 31263
rect 11713 31229 11747 31263
rect 11989 31229 12023 31263
rect 26249 31229 26283 31263
rect 27169 31229 27203 31263
rect 27629 31229 27663 31263
rect 11161 30889 11195 30923
rect 2881 30685 2915 30719
rect 11069 30685 11103 30719
rect 11897 30685 11931 30719
rect 14289 30685 14323 30719
rect 33977 30685 34011 30719
rect 2789 30209 2823 30243
rect 11805 30209 11839 30243
rect 14289 30209 14323 30243
rect 2973 30141 3007 30175
rect 4169 30141 4203 30175
rect 11989 30141 12023 30175
rect 12449 30141 12483 30175
rect 14473 30141 14507 30175
rect 14841 30141 14875 30175
rect 19441 30005 19475 30039
rect 27169 30005 27203 30039
rect 32965 30005 32999 30039
rect 33793 30005 33827 30039
rect 3157 29801 3191 29835
rect 12173 29801 12207 29835
rect 14473 29801 14507 29835
rect 19349 29665 19383 29699
rect 19809 29665 19843 29699
rect 25697 29665 25731 29699
rect 33057 29665 33091 29699
rect 34161 29665 34195 29699
rect 3249 29597 3283 29631
rect 12265 29597 12299 29631
rect 14381 29597 14415 29631
rect 25237 29597 25271 29631
rect 27721 29597 27755 29631
rect 28365 29597 28399 29631
rect 19533 29529 19567 29563
rect 25421 29529 25455 29563
rect 33977 29529 34011 29563
rect 27629 29461 27663 29495
rect 19809 29257 19843 29291
rect 27261 29189 27295 29223
rect 31217 29189 31251 29223
rect 34161 29189 34195 29223
rect 19901 29121 19935 29155
rect 26157 29121 26191 29155
rect 27077 29121 27111 29155
rect 29377 29121 29411 29155
rect 32321 29121 32355 29155
rect 28457 29053 28491 29087
rect 29561 29053 29595 29087
rect 32505 29053 32539 29087
rect 25513 28917 25547 28951
rect 24961 28713 24995 28747
rect 27905 28713 27939 28747
rect 25513 28577 25547 28611
rect 27353 28577 27387 28611
rect 33517 28577 33551 28611
rect 34161 28577 34195 28611
rect 24869 28509 24903 28543
rect 27813 28509 27847 28543
rect 25697 28441 25731 28475
rect 33977 28441 34011 28475
rect 25513 28169 25547 28203
rect 32781 28169 32815 28203
rect 33425 28169 33459 28203
rect 34069 28169 34103 28203
rect 25421 28033 25455 28067
rect 32873 28033 32907 28067
rect 33517 28033 33551 28067
rect 33977 28033 34011 28067
rect 31309 26741 31343 26775
rect 31309 26401 31343 26435
rect 33057 26401 33091 26435
rect 8125 26333 8159 26367
rect 29837 26333 29871 26367
rect 31493 26265 31527 26299
rect 32229 25993 32263 26027
rect 7849 25925 7883 25959
rect 31585 25925 31619 25959
rect 9689 25857 9723 25891
rect 29101 25857 29135 25891
rect 29745 25857 29779 25891
rect 32137 25857 32171 25891
rect 9505 25789 9539 25823
rect 29193 25789 29227 25823
rect 29929 25789 29963 25823
rect 10149 25653 10183 25687
rect 9045 25449 9079 25483
rect 9965 25313 9999 25347
rect 10425 25313 10459 25347
rect 32965 25313 32999 25347
rect 7757 25245 7791 25279
rect 9137 25245 9171 25279
rect 31033 25245 31067 25279
rect 31493 25245 31527 25279
rect 10149 25177 10183 25211
rect 31677 25177 31711 25211
rect 10333 24905 10367 24939
rect 31217 24905 31251 24939
rect 7665 24769 7699 24803
rect 10425 24769 10459 24803
rect 31125 24769 31159 24803
rect 7849 24701 7883 24735
rect 8401 24701 8435 24735
rect 32505 24565 32539 24599
rect 8309 24361 8343 24395
rect 8401 24157 8435 24191
rect 29837 24157 29871 24191
rect 30849 24157 30883 24191
rect 32137 24157 32171 24191
rect 32781 24157 32815 24191
rect 19717 24089 19751 24123
rect 19993 24021 20027 24055
rect 29929 24021 29963 24055
rect 32229 24021 32263 24055
rect 17509 23817 17543 23851
rect 18245 23749 18279 23783
rect 29929 23749 29963 23783
rect 32505 23749 32539 23783
rect 34161 23749 34195 23783
rect 17325 23681 17359 23715
rect 17969 23681 18003 23715
rect 19257 23681 19291 23715
rect 20177 23681 20211 23715
rect 32321 23681 32355 23715
rect 29745 23613 29779 23647
rect 30205 23613 30239 23647
rect 19349 23477 19383 23511
rect 20453 23477 20487 23511
rect 29837 23273 29871 23307
rect 30849 23137 30883 23171
rect 32689 23137 32723 23171
rect 19993 23069 20027 23103
rect 33149 23069 33183 23103
rect 31033 23001 31067 23035
rect 19717 22933 19751 22967
rect 33241 22933 33275 22967
rect 30849 22729 30883 22763
rect 32505 22661 32539 22695
rect 34161 22661 34195 22695
rect 30757 22593 30791 22627
rect 32321 22525 32355 22559
rect 17693 21505 17727 21539
rect 17509 21437 17543 21471
rect 17325 20893 17359 20927
rect 28365 20893 28399 20927
rect 29561 20893 29595 20927
rect 17601 20757 17635 20791
rect 30205 20485 30239 20519
rect 9229 20417 9263 20451
rect 15945 20417 15979 20451
rect 16957 20417 16991 20451
rect 17233 20417 17267 20451
rect 18705 20417 18739 20451
rect 27721 20417 27755 20451
rect 28365 20417 28399 20451
rect 18521 20349 18555 20383
rect 27813 20349 27847 20383
rect 28549 20349 28583 20383
rect 8585 20213 8619 20247
rect 9137 20213 9171 20247
rect 16129 20213 16163 20247
rect 24685 20213 24719 20247
rect 16313 20009 16347 20043
rect 11529 19873 11563 19907
rect 17049 19873 17083 19907
rect 24593 19873 24627 19907
rect 29561 19873 29595 19907
rect 9413 19805 9447 19839
rect 10609 19805 10643 19839
rect 11069 19805 11103 19839
rect 17325 19805 17359 19839
rect 28825 19805 28859 19839
rect 11253 19737 11287 19771
rect 16221 19737 16255 19771
rect 24777 19737 24811 19771
rect 26433 19737 26467 19771
rect 28917 19737 28951 19771
rect 29745 19737 29779 19771
rect 31401 19737 31435 19771
rect 11621 19465 11655 19499
rect 24317 19465 24351 19499
rect 8677 19397 8711 19431
rect 18061 19397 18095 19431
rect 18981 19397 19015 19431
rect 8493 19329 8527 19363
rect 10333 19329 10367 19363
rect 11713 19329 11747 19363
rect 16865 19329 16899 19363
rect 17785 19329 17819 19363
rect 18705 19329 18739 19363
rect 24225 19329 24259 19363
rect 17141 19261 17175 19295
rect 33057 19261 33091 19295
rect 33977 19261 34011 19295
rect 34161 19261 34195 19295
rect 6377 19125 6411 19159
rect 10793 19125 10827 19159
rect 17509 18921 17543 18955
rect 33241 18921 33275 18955
rect 33977 18921 34011 18955
rect 6285 18785 6319 18819
rect 10241 18785 10275 18819
rect 10701 18785 10735 18819
rect 29009 18785 29043 18819
rect 5273 18717 5307 18751
rect 9137 18717 9171 18751
rect 9597 18717 9631 18751
rect 16773 18717 16807 18751
rect 27169 18717 27203 18751
rect 31677 18717 31711 18751
rect 32321 18717 32355 18751
rect 33149 18717 33183 18751
rect 6469 18649 6503 18683
rect 8125 18649 8159 18683
rect 9689 18649 9723 18683
rect 10425 18649 10459 18683
rect 17417 18649 17451 18683
rect 18337 18649 18371 18683
rect 27353 18649 27387 18683
rect 9045 18581 9079 18615
rect 16497 18581 16531 18615
rect 18613 18581 18647 18615
rect 31769 18581 31803 18615
rect 6653 18377 6687 18411
rect 10977 18309 11011 18343
rect 18061 18309 18095 18343
rect 32321 18309 32355 18343
rect 6745 18241 6779 18275
rect 7849 18241 7883 18275
rect 9137 18241 9171 18275
rect 17417 18241 17451 18275
rect 27537 18241 27571 18275
rect 32137 18241 32171 18275
rect 9321 18173 9355 18207
rect 33885 18173 33919 18207
rect 7941 18037 7975 18071
rect 8677 18037 8711 18071
rect 17141 18037 17175 18071
rect 18337 18037 18371 18071
rect 29561 18037 29595 18071
rect 27261 17833 27295 17867
rect 5181 17697 5215 17731
rect 6837 17697 6871 17731
rect 8953 17697 8987 17731
rect 9413 17697 9447 17731
rect 29561 17697 29595 17731
rect 31401 17697 31435 17731
rect 2053 17629 2087 17663
rect 2789 17629 2823 17663
rect 17601 17629 17635 17663
rect 27169 17629 27203 17663
rect 27997 17629 28031 17663
rect 28825 17629 28859 17663
rect 5365 17561 5399 17595
rect 9137 17561 9171 17595
rect 28917 17561 28951 17595
rect 29745 17561 29779 17595
rect 1961 17493 1995 17527
rect 17509 17493 17543 17527
rect 27905 17493 27939 17527
rect 5365 17289 5399 17323
rect 27721 17221 27755 17255
rect 2329 17153 2363 17187
rect 2789 17153 2823 17187
rect 5273 17153 5307 17187
rect 2237 17085 2271 17119
rect 2973 17085 3007 17119
rect 3341 17085 3375 17119
rect 27537 17085 27571 17119
rect 29377 17085 29411 17119
rect 1501 16949 1535 16983
rect 32873 16949 32907 16983
rect 27629 16745 27663 16779
rect 1409 16609 1443 16643
rect 1593 16609 1627 16643
rect 32321 16609 32355 16643
rect 3249 16541 3283 16575
rect 32505 16473 32539 16507
rect 34161 16473 34195 16507
rect 32781 16201 32815 16235
rect 17417 16133 17451 16167
rect 9137 16065 9171 16099
rect 32873 16065 32907 16099
rect 21281 15997 21315 16031
rect 21833 15997 21867 16031
rect 22017 15997 22051 16031
rect 23673 15997 23707 16031
rect 4261 15861 4295 15895
rect 8493 15861 8527 15895
rect 9045 15861 9079 15895
rect 17141 15861 17175 15895
rect 20821 15657 20855 15691
rect 4261 15521 4295 15555
rect 4721 15521 4755 15555
rect 8953 15521 8987 15555
rect 9137 15521 9171 15555
rect 9873 15521 9907 15555
rect 17693 15453 17727 15487
rect 20729 15453 20763 15487
rect 4445 15385 4479 15419
rect 17509 15317 17543 15351
rect 4813 15113 4847 15147
rect 1961 14977 1995 15011
rect 4905 14977 4939 15011
rect 18889 14977 18923 15011
rect 25237 14977 25271 15011
rect 19165 14909 19199 14943
rect 1869 14773 1903 14807
rect 25329 14773 25363 14807
rect 1593 14433 1627 14467
rect 1869 14433 1903 14467
rect 25513 14433 25547 14467
rect 1409 14365 1443 14399
rect 25329 14365 25363 14399
rect 27169 14297 27203 14331
rect 1501 13889 1535 13923
rect 6561 13889 6595 13923
rect 17693 13889 17727 13923
rect 25329 13889 25363 13923
rect 5457 13821 5491 13855
rect 6469 13821 6503 13855
rect 16865 13685 16899 13719
rect 17601 13685 17635 13719
rect 25973 13685 26007 13719
rect 32781 13685 32815 13719
rect 33977 13685 34011 13719
rect 5273 13345 5307 13379
rect 7113 13345 7147 13379
rect 16865 13345 16899 13379
rect 17049 13345 17083 13379
rect 17325 13345 17359 13379
rect 25421 13345 25455 13379
rect 27261 13345 27295 13379
rect 33057 13345 33091 13379
rect 34161 13345 34195 13379
rect 7757 13277 7791 13311
rect 10241 13277 10275 13311
rect 6929 13209 6963 13243
rect 25605 13209 25639 13243
rect 33977 13209 34011 13243
rect 10425 13141 10459 13175
rect 25421 12937 25455 12971
rect 5733 12869 5767 12903
rect 8033 12869 8067 12903
rect 34161 12869 34195 12903
rect 5641 12801 5675 12835
rect 8217 12801 8251 12835
rect 25329 12801 25363 12835
rect 32321 12801 32355 12835
rect 6377 12733 6411 12767
rect 32505 12733 32539 12767
rect 32597 12393 32631 12427
rect 33885 12393 33919 12427
rect 32505 12189 32539 12223
rect 33793 12189 33827 12223
rect 17601 11713 17635 11747
rect 20729 11713 20763 11747
rect 14289 11509 14323 11543
rect 16957 11509 16991 11543
rect 17509 11509 17543 11543
rect 20821 11509 20855 11543
rect 14289 11169 14323 11203
rect 14841 11169 14875 11203
rect 16865 11169 16899 11203
rect 17049 11169 17083 11203
rect 17325 11169 17359 11203
rect 20913 11169 20947 11203
rect 21741 11169 21775 11203
rect 2329 11101 2363 11135
rect 2973 11101 3007 11135
rect 7297 11101 7331 11135
rect 9229 11101 9263 11135
rect 20729 11101 20763 11135
rect 5457 11033 5491 11067
rect 7113 11033 7147 11067
rect 14473 11033 14507 11067
rect 2881 10965 2915 10999
rect 6469 10761 6503 10795
rect 14473 10761 14507 10795
rect 2605 10693 2639 10727
rect 27261 10693 27295 10727
rect 27997 10693 28031 10727
rect 2421 10625 2455 10659
rect 6561 10625 6595 10659
rect 9137 10625 9171 10659
rect 14381 10625 14415 10659
rect 20729 10625 20763 10659
rect 27169 10625 27203 10659
rect 2881 10557 2915 10591
rect 5733 10557 5767 10591
rect 9321 10557 9355 10591
rect 9873 10557 9907 10591
rect 27813 10557 27847 10591
rect 29653 10557 29687 10591
rect 9781 10217 9815 10251
rect 27905 10217 27939 10251
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 9873 10013 9907 10047
rect 11345 10013 11379 10047
rect 11989 10013 12023 10047
rect 19533 10013 19567 10047
rect 1685 9877 1719 9911
rect 2973 9877 3007 9911
rect 11437 9877 11471 9911
rect 19625 9877 19659 9911
rect 2697 9605 2731 9639
rect 12081 9605 12115 9639
rect 19625 9605 19659 9639
rect 2513 9537 2547 9571
rect 11897 9537 11931 9571
rect 2973 9469 3007 9503
rect 13461 9469 13495 9503
rect 19441 9469 19475 9503
rect 19993 9469 20027 9503
rect 1501 9333 1535 9367
rect 19533 9129 19567 9163
rect 1409 8993 1443 9027
rect 1593 8993 1627 9027
rect 1869 8993 1903 9027
rect 23857 8925 23891 8959
rect 24593 8925 24627 8959
rect 30941 8925 30975 8959
rect 31125 8857 31159 8891
rect 32781 8857 32815 8891
rect 24501 8789 24535 8823
rect 30849 8585 30883 8619
rect 24133 8517 24167 8551
rect 11713 8449 11747 8483
rect 23949 8449 23983 8483
rect 29101 8449 29135 8483
rect 30757 8449 30791 8483
rect 31401 8449 31435 8483
rect 11621 8381 11655 8415
rect 24501 8381 24535 8415
rect 12357 8313 12391 8347
rect 29193 8245 29227 8279
rect 29745 8245 29779 8279
rect 12909 7905 12943 7939
rect 13093 7905 13127 7939
rect 29561 7905 29595 7939
rect 2421 7837 2455 7871
rect 11253 7769 11287 7803
rect 29745 7769 29779 7803
rect 31401 7769 31435 7803
rect 2421 7361 2455 7395
rect 6653 7361 6687 7395
rect 20729 7361 20763 7395
rect 2605 7293 2639 7327
rect 3157 7293 3191 7327
rect 6561 7157 6595 7191
rect 7297 7157 7331 7191
rect 20085 7157 20119 7191
rect 20821 7157 20855 7191
rect 32689 7157 32723 7191
rect 2973 6817 3007 6851
rect 8033 6817 8067 6851
rect 20085 6817 20119 6851
rect 20269 6817 20303 6851
rect 21465 6817 21499 6851
rect 32321 6817 32355 6851
rect 34161 6817 34195 6851
rect 3065 6749 3099 6783
rect 9781 6749 9815 6783
rect 10241 6749 10275 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 14105 6749 14139 6783
rect 27261 6749 27295 6783
rect 30573 6749 30607 6783
rect 31217 6749 31251 6783
rect 6193 6681 6227 6715
rect 7849 6681 7883 6715
rect 32505 6681 32539 6715
rect 9689 6613 9723 6647
rect 13369 6613 13403 6647
rect 14197 6613 14231 6647
rect 30665 6613 30699 6647
rect 32597 6409 32631 6443
rect 13001 6341 13035 6375
rect 10701 6273 10735 6307
rect 12817 6273 12851 6307
rect 27261 6273 27295 6307
rect 32505 6273 32539 6307
rect 7481 6205 7515 6239
rect 7941 6205 7975 6239
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 13277 6205 13311 6239
rect 27445 6205 27479 6239
rect 29101 6205 29135 6239
rect 10609 6069 10643 6103
rect 15301 6069 15335 6103
rect 26985 5865 27019 5899
rect 6561 5729 6595 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 10609 5729 10643 5763
rect 15761 5729 15795 5763
rect 15945 5729 15979 5763
rect 30665 5729 30699 5763
rect 30849 5729 30883 5763
rect 32229 5729 32263 5763
rect 9137 5661 9171 5695
rect 26893 5661 26927 5695
rect 27629 5661 27663 5695
rect 6745 5593 6779 5627
rect 8401 5593 8435 5627
rect 14105 5593 14139 5627
rect 7849 5321 7883 5355
rect 9229 5253 9263 5287
rect 7113 5185 7147 5219
rect 7941 5185 7975 5219
rect 9045 5185 9079 5219
rect 11713 5185 11747 5219
rect 27537 5185 27571 5219
rect 30297 5185 30331 5219
rect 10793 5117 10827 5151
rect 27721 5117 27755 5151
rect 29377 5117 29411 5151
rect 6653 4981 6687 5015
rect 8585 4981 8619 5015
rect 11621 4981 11655 5015
rect 30389 4981 30423 5015
rect 7941 4777 7975 4811
rect 27353 4777 27387 4811
rect 10977 4641 11011 4675
rect 11161 4641 11195 4675
rect 30481 4641 30515 4675
rect 30941 4641 30975 4675
rect 7389 4573 7423 4607
rect 8033 4573 8067 4607
rect 27261 4573 27295 4607
rect 30297 4573 30331 4607
rect 9321 4505 9355 4539
rect 7297 4437 7331 4471
rect 7297 4165 7331 4199
rect 7113 4097 7147 4131
rect 9873 4097 9907 4131
rect 30297 4097 30331 4131
rect 32229 4097 32263 4131
rect 7573 4029 7607 4063
rect 9965 3893 9999 3927
rect 10517 3893 10551 3927
rect 32321 3893 32355 3927
rect 32873 3893 32907 3927
rect 9781 3553 9815 3587
rect 9965 3553 9999 3587
rect 10333 3553 10367 3587
rect 16129 3553 16163 3587
rect 32321 3553 32355 3587
rect 32505 3553 32539 3587
rect 2789 3485 2823 3519
rect 15577 3485 15611 3519
rect 17877 3485 17911 3519
rect 15761 3417 15795 3451
rect 34161 3417 34195 3451
rect 17049 3077 17083 3111
rect 17785 3077 17819 3111
rect 2789 3009 2823 3043
rect 15577 3009 15611 3043
rect 16957 3009 16991 3043
rect 17601 3009 17635 3043
rect 2973 2941 3007 2975
rect 3249 2941 3283 2975
rect 19441 2941 19475 2975
rect 3157 2601 3191 2635
rect 15761 2601 15795 2635
rect 3249 2397 3283 2431
rect 15669 2397 15703 2431
<< metal1 >>
rect 29730 40060 29736 40112
rect 29788 40100 29794 40112
rect 31754 40100 31760 40112
rect 29788 40072 31760 40100
rect 29788 40060 29794 40072
rect 31754 40060 31760 40072
rect 31812 40060 31818 40112
rect 1104 39738 34868 39760
rect 1104 39686 5174 39738
rect 5226 39686 5238 39738
rect 5290 39686 5302 39738
rect 5354 39686 5366 39738
rect 5418 39686 5430 39738
rect 5482 39686 13622 39738
rect 13674 39686 13686 39738
rect 13738 39686 13750 39738
rect 13802 39686 13814 39738
rect 13866 39686 13878 39738
rect 13930 39686 22070 39738
rect 22122 39686 22134 39738
rect 22186 39686 22198 39738
rect 22250 39686 22262 39738
rect 22314 39686 22326 39738
rect 22378 39686 30518 39738
rect 30570 39686 30582 39738
rect 30634 39686 30646 39738
rect 30698 39686 30710 39738
rect 30762 39686 30774 39738
rect 30826 39686 34868 39738
rect 1104 39664 34868 39686
rect 17052 39460 19564 39488
rect 17052 39432 17080 39460
rect 7834 39420 7840 39432
rect 7795 39392 7840 39420
rect 7834 39380 7840 39392
rect 7892 39380 7898 39432
rect 16114 39420 16120 39432
rect 16075 39392 16120 39420
rect 16114 39380 16120 39392
rect 16172 39380 16178 39432
rect 17034 39420 17040 39432
rect 16995 39392 17040 39420
rect 17034 39380 17040 39392
rect 17092 39380 17098 39432
rect 19536 39429 19564 39460
rect 17681 39423 17739 39429
rect 17681 39389 17693 39423
rect 17727 39389 17739 39423
rect 17681 39383 17739 39389
rect 19521 39423 19579 39429
rect 19521 39389 19533 39423
rect 19567 39389 19579 39423
rect 19521 39383 19579 39389
rect 20349 39423 20407 39429
rect 20349 39389 20361 39423
rect 20395 39389 20407 39423
rect 20990 39420 20996 39432
rect 20951 39392 20996 39420
rect 20349 39383 20407 39389
rect 16942 39312 16948 39364
rect 17000 39352 17006 39364
rect 17696 39352 17724 39383
rect 17000 39324 17724 39352
rect 20364 39352 20392 39383
rect 20990 39380 20996 39392
rect 21048 39380 21054 39432
rect 22370 39380 22376 39432
rect 22428 39420 22434 39432
rect 22465 39423 22523 39429
rect 22465 39420 22477 39423
rect 22428 39392 22477 39420
rect 22428 39380 22434 39392
rect 22465 39389 22477 39392
rect 22511 39389 22523 39423
rect 22465 39383 22523 39389
rect 21082 39352 21088 39364
rect 20364 39324 21088 39352
rect 17000 39312 17006 39324
rect 21082 39312 21088 39324
rect 21140 39312 21146 39364
rect 17126 39284 17132 39296
rect 17087 39256 17132 39284
rect 17126 39244 17132 39256
rect 17184 39244 17190 39296
rect 18046 39244 18052 39296
rect 18104 39284 18110 39296
rect 19242 39284 19248 39296
rect 18104 39256 19248 39284
rect 18104 39244 18110 39256
rect 19242 39244 19248 39256
rect 19300 39244 19306 39296
rect 19613 39287 19671 39293
rect 19613 39253 19625 39287
rect 19659 39284 19671 39287
rect 20806 39284 20812 39296
rect 19659 39256 20812 39284
rect 19659 39253 19671 39256
rect 19613 39247 19671 39253
rect 20806 39244 20812 39256
rect 20864 39244 20870 39296
rect 1104 39194 34868 39216
rect 1104 39142 9398 39194
rect 9450 39142 9462 39194
rect 9514 39142 9526 39194
rect 9578 39142 9590 39194
rect 9642 39142 9654 39194
rect 9706 39142 17846 39194
rect 17898 39142 17910 39194
rect 17962 39142 17974 39194
rect 18026 39142 18038 39194
rect 18090 39142 18102 39194
rect 18154 39142 26294 39194
rect 26346 39142 26358 39194
rect 26410 39142 26422 39194
rect 26474 39142 26486 39194
rect 26538 39142 26550 39194
rect 26602 39142 34868 39194
rect 1104 39120 34868 39142
rect 17126 39012 17132 39024
rect 17087 38984 17132 39012
rect 17126 38972 17132 38984
rect 17184 38972 17190 39024
rect 24213 39015 24271 39021
rect 24213 38981 24225 39015
rect 24259 39012 24271 39015
rect 25130 39012 25136 39024
rect 24259 38984 25136 39012
rect 24259 38981 24271 38984
rect 24213 38975 24271 38981
rect 25130 38972 25136 38984
rect 25188 38972 25194 39024
rect 7834 38944 7840 38956
rect 7795 38916 7840 38944
rect 7834 38904 7840 38916
rect 7892 38904 7898 38956
rect 16117 38947 16175 38953
rect 16117 38913 16129 38947
rect 16163 38944 16175 38947
rect 16942 38944 16948 38956
rect 16163 38916 16574 38944
rect 16903 38916 16948 38944
rect 16163 38913 16175 38916
rect 16117 38907 16175 38913
rect 8018 38876 8024 38888
rect 7979 38848 8024 38876
rect 8018 38836 8024 38848
rect 8076 38836 8082 38888
rect 8386 38876 8392 38888
rect 8347 38848 8392 38876
rect 8386 38836 8392 38848
rect 8444 38836 8450 38888
rect 16546 38808 16574 38916
rect 16942 38904 16948 38916
rect 17000 38904 17006 38956
rect 21082 38904 21088 38956
rect 21140 38944 21146 38956
rect 22370 38944 22376 38956
rect 21140 38916 21185 38944
rect 22331 38916 22376 38944
rect 21140 38904 21146 38916
rect 22370 38904 22376 38916
rect 22428 38904 22434 38956
rect 17402 38876 17408 38888
rect 17363 38848 17408 38876
rect 17402 38836 17408 38848
rect 17460 38836 17466 38888
rect 19334 38876 19340 38888
rect 19295 38848 19340 38876
rect 19334 38836 19340 38848
rect 19392 38836 19398 38888
rect 20898 38876 20904 38888
rect 20859 38848 20904 38876
rect 20898 38836 20904 38848
rect 20956 38836 20962 38888
rect 22554 38876 22560 38888
rect 22515 38848 22560 38876
rect 22554 38836 22560 38848
rect 22612 38836 22618 38888
rect 17034 38808 17040 38820
rect 16546 38780 17040 38808
rect 17034 38768 17040 38780
rect 17092 38768 17098 38820
rect 20254 38768 20260 38820
rect 20312 38808 20318 38820
rect 31754 38808 31760 38820
rect 20312 38780 31760 38808
rect 20312 38768 20318 38780
rect 31754 38768 31760 38780
rect 31812 38768 31818 38820
rect 4890 38700 4896 38752
rect 4948 38740 4954 38752
rect 4985 38743 5043 38749
rect 4985 38740 4997 38743
rect 4948 38712 4997 38740
rect 4948 38700 4954 38712
rect 4985 38709 4997 38712
rect 5031 38709 5043 38743
rect 4985 38703 5043 38709
rect 16025 38743 16083 38749
rect 16025 38709 16037 38743
rect 16071 38740 16083 38743
rect 16574 38740 16580 38752
rect 16071 38712 16580 38740
rect 16071 38709 16083 38712
rect 16025 38703 16083 38709
rect 16574 38700 16580 38712
rect 16632 38700 16638 38752
rect 28442 38700 28448 38752
rect 28500 38740 28506 38752
rect 28537 38743 28595 38749
rect 28537 38740 28549 38743
rect 28500 38712 28549 38740
rect 28500 38700 28506 38712
rect 28537 38709 28549 38712
rect 28583 38709 28595 38743
rect 28537 38703 28595 38709
rect 1104 38650 34868 38672
rect 1104 38598 5174 38650
rect 5226 38598 5238 38650
rect 5290 38598 5302 38650
rect 5354 38598 5366 38650
rect 5418 38598 5430 38650
rect 5482 38598 13622 38650
rect 13674 38598 13686 38650
rect 13738 38598 13750 38650
rect 13802 38598 13814 38650
rect 13866 38598 13878 38650
rect 13930 38598 22070 38650
rect 22122 38598 22134 38650
rect 22186 38598 22198 38650
rect 22250 38598 22262 38650
rect 22314 38598 22326 38650
rect 22378 38598 30518 38650
rect 30570 38598 30582 38650
rect 30634 38598 30646 38650
rect 30698 38598 30710 38650
rect 30762 38598 30774 38650
rect 30826 38598 34868 38650
rect 1104 38576 34868 38598
rect 14 38496 20 38548
rect 72 38536 78 38548
rect 1302 38536 1308 38548
rect 72 38508 1308 38536
rect 72 38496 78 38508
rect 1302 38496 1308 38508
rect 1360 38496 1366 38548
rect 8018 38536 8024 38548
rect 7979 38508 8024 38536
rect 8018 38496 8024 38508
rect 8076 38496 8082 38548
rect 22373 38539 22431 38545
rect 22373 38505 22385 38539
rect 22419 38536 22431 38539
rect 22554 38536 22560 38548
rect 22419 38508 22560 38536
rect 22419 38505 22431 38508
rect 22373 38499 22431 38505
rect 22554 38496 22560 38508
rect 22612 38496 22618 38548
rect 4062 38428 4068 38480
rect 4120 38468 4126 38480
rect 4120 38440 5580 38468
rect 4120 38428 4126 38440
rect 4890 38400 4896 38412
rect 4851 38372 4896 38400
rect 4890 38360 4896 38372
rect 4948 38360 4954 38412
rect 5552 38409 5580 38440
rect 9030 38428 9036 38480
rect 9088 38468 9094 38480
rect 19334 38468 19340 38480
rect 9088 38440 19340 38468
rect 9088 38428 9094 38440
rect 19334 38428 19340 38440
rect 19392 38428 19398 38480
rect 19978 38428 19984 38480
rect 20036 38428 20042 38480
rect 5537 38403 5595 38409
rect 5537 38369 5549 38403
rect 5583 38369 5595 38403
rect 5537 38363 5595 38369
rect 16114 38360 16120 38412
rect 16172 38400 16178 38412
rect 16393 38403 16451 38409
rect 16393 38400 16405 38403
rect 16172 38372 16405 38400
rect 16172 38360 16178 38372
rect 16393 38369 16405 38372
rect 16439 38369 16451 38403
rect 16393 38363 16451 38369
rect 16574 38360 16580 38412
rect 16632 38400 16638 38412
rect 16850 38400 16856 38412
rect 16632 38372 16677 38400
rect 16811 38372 16856 38400
rect 16632 38360 16638 38372
rect 16850 38360 16856 38372
rect 16908 38360 16914 38412
rect 19889 38403 19947 38409
rect 19889 38369 19901 38403
rect 19935 38400 19947 38403
rect 19996 38400 20024 38428
rect 19935 38372 20024 38400
rect 19935 38369 19947 38372
rect 19889 38363 19947 38369
rect 20990 38360 20996 38412
rect 21048 38400 21054 38412
rect 21269 38403 21327 38409
rect 21269 38400 21281 38403
rect 21048 38372 21281 38400
rect 21048 38360 21054 38372
rect 21269 38369 21281 38372
rect 21315 38369 21327 38403
rect 21269 38363 21327 38369
rect 6730 38292 6736 38344
rect 6788 38332 6794 38344
rect 7929 38335 7987 38341
rect 7929 38332 7941 38335
rect 6788 38304 7941 38332
rect 6788 38292 6794 38304
rect 7929 38301 7941 38304
rect 7975 38301 7987 38335
rect 7929 38295 7987 38301
rect 22281 38335 22339 38341
rect 22281 38301 22293 38335
rect 22327 38332 22339 38335
rect 23474 38332 23480 38344
rect 22327 38304 23480 38332
rect 22327 38301 22339 38304
rect 22281 38295 22339 38301
rect 23474 38292 23480 38304
rect 23532 38292 23538 38344
rect 28258 38292 28264 38344
rect 28316 38332 28322 38344
rect 28537 38335 28595 38341
rect 28537 38332 28549 38335
rect 28316 38304 28549 38332
rect 28316 38292 28322 38304
rect 28537 38301 28549 38304
rect 28583 38332 28595 38335
rect 30282 38332 30288 38344
rect 28583 38304 30288 38332
rect 28583 38301 28595 38304
rect 28537 38295 28595 38301
rect 30282 38292 30288 38304
rect 30340 38292 30346 38344
rect 32306 38292 32312 38344
rect 32364 38332 32370 38344
rect 32769 38335 32827 38341
rect 32769 38332 32781 38335
rect 32364 38304 32781 38332
rect 32364 38292 32370 38304
rect 32769 38301 32781 38304
rect 32815 38301 32827 38335
rect 32769 38295 32827 38301
rect 5077 38267 5135 38273
rect 5077 38233 5089 38267
rect 5123 38264 5135 38267
rect 5534 38264 5540 38276
rect 5123 38236 5540 38264
rect 5123 38233 5135 38236
rect 5077 38227 5135 38233
rect 5534 38224 5540 38236
rect 5592 38224 5598 38276
rect 20806 38224 20812 38276
rect 20864 38264 20870 38276
rect 21085 38267 21143 38273
rect 21085 38264 21097 38267
rect 20864 38236 21097 38264
rect 20864 38224 20870 38236
rect 21085 38233 21097 38236
rect 21131 38233 21143 38267
rect 21085 38227 21143 38233
rect 16206 38156 16212 38208
rect 16264 38196 16270 38208
rect 16850 38196 16856 38208
rect 16264 38168 16856 38196
rect 16264 38156 16270 38168
rect 16850 38156 16856 38168
rect 16908 38156 16914 38208
rect 28626 38196 28632 38208
rect 28587 38168 28632 38196
rect 28626 38156 28632 38168
rect 28684 38156 28690 38208
rect 1104 38106 34868 38128
rect 1104 38054 9398 38106
rect 9450 38054 9462 38106
rect 9514 38054 9526 38106
rect 9578 38054 9590 38106
rect 9642 38054 9654 38106
rect 9706 38054 17846 38106
rect 17898 38054 17910 38106
rect 17962 38054 17974 38106
rect 18026 38054 18038 38106
rect 18090 38054 18102 38106
rect 18154 38054 26294 38106
rect 26346 38054 26358 38106
rect 26410 38054 26422 38106
rect 26474 38054 26486 38106
rect 26538 38054 26550 38106
rect 26602 38054 34868 38106
rect 1104 38032 34868 38054
rect 5534 37992 5540 38004
rect 5495 37964 5540 37992
rect 5534 37952 5540 37964
rect 5592 37952 5598 38004
rect 19797 37995 19855 38001
rect 19797 37961 19809 37995
rect 19843 37992 19855 37995
rect 20898 37992 20904 38004
rect 19843 37964 20904 37992
rect 19843 37961 19855 37964
rect 19797 37955 19855 37961
rect 20898 37952 20904 37964
rect 20956 37952 20962 38004
rect 34054 37992 34060 38004
rect 26206 37964 34060 37992
rect 20070 37884 20076 37936
rect 20128 37924 20134 37936
rect 26206 37924 26234 37964
rect 34054 37952 34060 37964
rect 34112 37952 34118 38004
rect 28626 37924 28632 37936
rect 20128 37896 26234 37924
rect 28587 37896 28632 37924
rect 20128 37884 20134 37896
rect 28626 37884 28632 37896
rect 28684 37884 28690 37936
rect 34146 37924 34152 37936
rect 34107 37896 34152 37924
rect 34146 37884 34152 37896
rect 34204 37884 34210 37936
rect 5629 37859 5687 37865
rect 5629 37825 5641 37859
rect 5675 37856 5687 37859
rect 6730 37856 6736 37868
rect 5675 37828 6736 37856
rect 5675 37825 5687 37828
rect 5629 37819 5687 37825
rect 6730 37816 6736 37828
rect 6788 37816 6794 37868
rect 7098 37816 7104 37868
rect 7156 37856 7162 37868
rect 10410 37856 10416 37868
rect 7156 37828 10416 37856
rect 7156 37816 7162 37828
rect 10410 37816 10416 37828
rect 10468 37816 10474 37868
rect 19889 37859 19947 37865
rect 19889 37825 19901 37859
rect 19935 37856 19947 37859
rect 28258 37856 28264 37868
rect 19935 37828 28264 37856
rect 19935 37825 19947 37828
rect 19889 37819 19947 37825
rect 28258 37816 28264 37828
rect 28316 37816 28322 37868
rect 28442 37856 28448 37868
rect 28403 37828 28448 37856
rect 28442 37816 28448 37828
rect 28500 37816 28506 37868
rect 32306 37856 32312 37868
rect 32267 37828 32312 37856
rect 32306 37816 32312 37828
rect 32364 37816 32370 37868
rect 28994 37788 29000 37800
rect 28955 37760 29000 37788
rect 28994 37748 29000 37760
rect 29052 37748 29058 37800
rect 32490 37788 32496 37800
rect 32451 37760 32496 37788
rect 32490 37748 32496 37760
rect 32548 37748 32554 37800
rect 7285 37655 7343 37661
rect 7285 37621 7297 37655
rect 7331 37652 7343 37655
rect 8386 37652 8392 37664
rect 7331 37624 8392 37652
rect 7331 37621 7343 37624
rect 7285 37615 7343 37621
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 22097 37655 22155 37661
rect 22097 37621 22109 37655
rect 22143 37652 22155 37655
rect 22462 37652 22468 37664
rect 22143 37624 22468 37652
rect 22143 37621 22155 37624
rect 22097 37615 22155 37621
rect 22462 37612 22468 37624
rect 22520 37612 22526 37664
rect 1104 37562 34868 37584
rect 1104 37510 5174 37562
rect 5226 37510 5238 37562
rect 5290 37510 5302 37562
rect 5354 37510 5366 37562
rect 5418 37510 5430 37562
rect 5482 37510 13622 37562
rect 13674 37510 13686 37562
rect 13738 37510 13750 37562
rect 13802 37510 13814 37562
rect 13866 37510 13878 37562
rect 13930 37510 22070 37562
rect 22122 37510 22134 37562
rect 22186 37510 22198 37562
rect 22250 37510 22262 37562
rect 22314 37510 22326 37562
rect 22378 37510 30518 37562
rect 30570 37510 30582 37562
rect 30634 37510 30646 37562
rect 30698 37510 30710 37562
rect 30762 37510 30774 37562
rect 30826 37510 34868 37562
rect 1104 37488 34868 37510
rect 32490 37448 32496 37460
rect 32451 37420 32496 37448
rect 32490 37408 32496 37420
rect 32548 37408 32554 37460
rect 22462 37312 22468 37324
rect 22020 37284 22468 37312
rect 658 37204 664 37256
rect 716 37244 722 37256
rect 6549 37247 6607 37253
rect 6549 37244 6561 37247
rect 716 37216 6561 37244
rect 716 37204 722 37216
rect 6549 37213 6561 37216
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 8444 37216 8489 37244
rect 8444 37204 8450 37216
rect 18414 37204 18420 37256
rect 18472 37244 18478 37256
rect 22020 37253 22048 37284
rect 22462 37272 22468 37284
rect 22520 37272 22526 37324
rect 22646 37312 22652 37324
rect 22607 37284 22652 37312
rect 22646 37272 22652 37284
rect 22704 37272 22710 37324
rect 30282 37272 30288 37324
rect 30340 37312 30346 37324
rect 30340 37284 32444 37312
rect 30340 37272 30346 37284
rect 32416 37253 32444 37284
rect 18509 37247 18567 37253
rect 18509 37244 18521 37247
rect 18472 37216 18521 37244
rect 18472 37204 18478 37216
rect 18509 37213 18521 37216
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 22005 37247 22063 37253
rect 22005 37213 22017 37247
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 32401 37247 32459 37253
rect 32401 37213 32413 37247
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 7374 37136 7380 37188
rect 7432 37176 7438 37188
rect 8205 37179 8263 37185
rect 8205 37176 8217 37179
rect 7432 37148 8217 37176
rect 7432 37136 7438 37148
rect 8205 37145 8217 37148
rect 8251 37145 8263 37179
rect 22186 37176 22192 37188
rect 22147 37148 22192 37176
rect 8205 37139 8263 37145
rect 22186 37136 22192 37148
rect 22244 37136 22250 37188
rect 1104 37018 34868 37040
rect 1104 36966 9398 37018
rect 9450 36966 9462 37018
rect 9514 36966 9526 37018
rect 9578 36966 9590 37018
rect 9642 36966 9654 37018
rect 9706 36966 17846 37018
rect 17898 36966 17910 37018
rect 17962 36966 17974 37018
rect 18026 36966 18038 37018
rect 18090 36966 18102 37018
rect 18154 36966 26294 37018
rect 26346 36966 26358 37018
rect 26410 36966 26422 37018
rect 26474 36966 26486 37018
rect 26538 36966 26550 37018
rect 26602 36966 34868 37018
rect 1104 36944 34868 36966
rect 7374 36904 7380 36916
rect 7335 36876 7380 36904
rect 7374 36864 7380 36876
rect 7432 36864 7438 36916
rect 22186 36904 22192 36916
rect 22147 36876 22192 36904
rect 22186 36864 22192 36876
rect 22244 36864 22250 36916
rect 20254 36836 20260 36848
rect 20215 36808 20260 36836
rect 20254 36796 20260 36808
rect 20312 36796 20318 36848
rect 7469 36771 7527 36777
rect 7469 36737 7481 36771
rect 7515 36768 7527 36771
rect 17494 36768 17500 36780
rect 7515 36740 17500 36768
rect 7515 36737 7527 36740
rect 7469 36731 7527 36737
rect 17494 36728 17500 36740
rect 17552 36768 17558 36780
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17552 36740 17785 36768
rect 17552 36728 17558 36740
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 18414 36768 18420 36780
rect 18375 36740 18420 36768
rect 17773 36731 17831 36737
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 22097 36771 22155 36777
rect 22097 36737 22109 36771
rect 22143 36768 22155 36771
rect 27798 36768 27804 36780
rect 22143 36740 27804 36768
rect 22143 36737 22155 36740
rect 22097 36731 22155 36737
rect 27798 36728 27804 36740
rect 27856 36728 27862 36780
rect 17865 36703 17923 36709
rect 17865 36669 17877 36703
rect 17911 36700 17923 36703
rect 18601 36703 18659 36709
rect 18601 36700 18613 36703
rect 17911 36672 18613 36700
rect 17911 36669 17923 36672
rect 17865 36663 17923 36669
rect 18601 36669 18613 36672
rect 18647 36669 18659 36703
rect 18601 36663 18659 36669
rect 17310 36564 17316 36576
rect 17271 36536 17316 36564
rect 17310 36524 17316 36536
rect 17368 36524 17374 36576
rect 1104 36474 34868 36496
rect 1104 36422 5174 36474
rect 5226 36422 5238 36474
rect 5290 36422 5302 36474
rect 5354 36422 5366 36474
rect 5418 36422 5430 36474
rect 5482 36422 13622 36474
rect 13674 36422 13686 36474
rect 13738 36422 13750 36474
rect 13802 36422 13814 36474
rect 13866 36422 13878 36474
rect 13930 36422 22070 36474
rect 22122 36422 22134 36474
rect 22186 36422 22198 36474
rect 22250 36422 22262 36474
rect 22314 36422 22326 36474
rect 22378 36422 30518 36474
rect 30570 36422 30582 36474
rect 30634 36422 30646 36474
rect 30698 36422 30710 36474
rect 30762 36422 30774 36474
rect 30826 36422 34868 36474
rect 1104 36400 34868 36422
rect 17494 36156 17500 36168
rect 17455 36128 17500 36156
rect 17494 36116 17500 36128
rect 17552 36116 17558 36168
rect 27890 36156 27896 36168
rect 27851 36128 27896 36156
rect 27890 36116 27896 36128
rect 27948 36116 27954 36168
rect 1854 36088 1860 36100
rect 1815 36060 1860 36088
rect 1854 36048 1860 36060
rect 1912 36048 1918 36100
rect 1946 36020 1952 36032
rect 1907 35992 1952 36020
rect 1946 35980 1952 35992
rect 2004 35980 2010 36032
rect 17589 36023 17647 36029
rect 17589 35989 17601 36023
rect 17635 36020 17647 36023
rect 17678 36020 17684 36032
rect 17635 35992 17684 36020
rect 17635 35989 17647 35992
rect 17589 35983 17647 35989
rect 17678 35980 17684 35992
rect 17736 35980 17742 36032
rect 1104 35930 34868 35952
rect 1104 35878 9398 35930
rect 9450 35878 9462 35930
rect 9514 35878 9526 35930
rect 9578 35878 9590 35930
rect 9642 35878 9654 35930
rect 9706 35878 17846 35930
rect 17898 35878 17910 35930
rect 17962 35878 17974 35930
rect 18026 35878 18038 35930
rect 18090 35878 18102 35930
rect 18154 35878 26294 35930
rect 26346 35878 26358 35930
rect 26410 35878 26422 35930
rect 26474 35878 26486 35930
rect 26538 35878 26550 35930
rect 26602 35878 34868 35930
rect 1104 35856 34868 35878
rect 17678 35748 17684 35760
rect 17639 35720 17684 35748
rect 17678 35708 17684 35720
rect 17736 35708 17742 35760
rect 29730 35748 29736 35760
rect 29691 35720 29736 35748
rect 29730 35708 29736 35720
rect 29788 35708 29794 35760
rect 17310 35640 17316 35692
rect 17368 35680 17374 35692
rect 17497 35683 17555 35689
rect 17497 35680 17509 35683
rect 17368 35652 17509 35680
rect 17368 35640 17374 35652
rect 17497 35649 17509 35652
rect 17543 35649 17555 35683
rect 27890 35680 27896 35692
rect 27851 35652 27896 35680
rect 17497 35643 17555 35649
rect 27890 35640 27896 35652
rect 27948 35640 27954 35692
rect 19242 35612 19248 35624
rect 19203 35584 19248 35612
rect 19242 35572 19248 35584
rect 19300 35572 19306 35624
rect 28074 35612 28080 35624
rect 28035 35584 28080 35612
rect 28074 35572 28080 35584
rect 28132 35572 28138 35624
rect 1104 35386 34868 35408
rect 1104 35334 5174 35386
rect 5226 35334 5238 35386
rect 5290 35334 5302 35386
rect 5354 35334 5366 35386
rect 5418 35334 5430 35386
rect 5482 35334 13622 35386
rect 13674 35334 13686 35386
rect 13738 35334 13750 35386
rect 13802 35334 13814 35386
rect 13866 35334 13878 35386
rect 13930 35334 22070 35386
rect 22122 35334 22134 35386
rect 22186 35334 22198 35386
rect 22250 35334 22262 35386
rect 22314 35334 22326 35386
rect 22378 35334 30518 35386
rect 30570 35334 30582 35386
rect 30634 35334 30646 35386
rect 30698 35334 30710 35386
rect 30762 35334 30774 35386
rect 30826 35334 34868 35386
rect 1104 35312 34868 35334
rect 27893 35275 27951 35281
rect 27893 35241 27905 35275
rect 27939 35272 27951 35275
rect 28074 35272 28080 35284
rect 27939 35244 28080 35272
rect 27939 35241 27951 35244
rect 27893 35235 27951 35241
rect 28074 35232 28080 35244
rect 28132 35232 28138 35284
rect 27798 35068 27804 35080
rect 27711 35040 27804 35068
rect 27798 35028 27804 35040
rect 27856 35068 27862 35080
rect 29086 35068 29092 35080
rect 27856 35040 29092 35068
rect 27856 35028 27862 35040
rect 29086 35028 29092 35040
rect 29144 35028 29150 35080
rect 1104 34842 34868 34864
rect 1104 34790 9398 34842
rect 9450 34790 9462 34842
rect 9514 34790 9526 34842
rect 9578 34790 9590 34842
rect 9642 34790 9654 34842
rect 9706 34790 17846 34842
rect 17898 34790 17910 34842
rect 17962 34790 17974 34842
rect 18026 34790 18038 34842
rect 18090 34790 18102 34842
rect 18154 34790 26294 34842
rect 26346 34790 26358 34842
rect 26410 34790 26422 34842
rect 26474 34790 26486 34842
rect 26538 34790 26550 34842
rect 26602 34790 34868 34842
rect 1104 34768 34868 34790
rect 9858 34348 9864 34400
rect 9916 34388 9922 34400
rect 9953 34391 10011 34397
rect 9953 34388 9965 34391
rect 9916 34360 9965 34388
rect 9916 34348 9922 34360
rect 9953 34357 9965 34360
rect 9999 34357 10011 34391
rect 9953 34351 10011 34357
rect 1104 34298 34868 34320
rect 1104 34246 5174 34298
rect 5226 34246 5238 34298
rect 5290 34246 5302 34298
rect 5354 34246 5366 34298
rect 5418 34246 5430 34298
rect 5482 34246 13622 34298
rect 13674 34246 13686 34298
rect 13738 34246 13750 34298
rect 13802 34246 13814 34298
rect 13866 34246 13878 34298
rect 13930 34246 22070 34298
rect 22122 34246 22134 34298
rect 22186 34246 22198 34298
rect 22250 34246 22262 34298
rect 22314 34246 22326 34298
rect 22378 34246 30518 34298
rect 30570 34246 30582 34298
rect 30634 34246 30646 34298
rect 30698 34246 30710 34298
rect 30762 34246 30774 34298
rect 30826 34246 34868 34298
rect 1104 34224 34868 34246
rect 6886 34088 10364 34116
rect 3418 33872 3424 33924
rect 3476 33912 3482 33924
rect 6886 33912 6914 34088
rect 9858 34048 9864 34060
rect 9819 34020 9864 34048
rect 9858 34008 9864 34020
rect 9916 34008 9922 34060
rect 10336 34057 10364 34088
rect 10321 34051 10379 34057
rect 10321 34017 10333 34051
rect 10367 34017 10379 34051
rect 10321 34011 10379 34017
rect 27614 33980 27620 33992
rect 27575 33952 27620 33980
rect 27614 33940 27620 33952
rect 27672 33940 27678 33992
rect 3476 33884 6914 33912
rect 10045 33915 10103 33921
rect 3476 33872 3482 33884
rect 10045 33881 10057 33915
rect 10091 33912 10103 33915
rect 10226 33912 10232 33924
rect 10091 33884 10232 33912
rect 10091 33881 10103 33884
rect 10045 33875 10103 33881
rect 10226 33872 10232 33884
rect 10284 33872 10290 33924
rect 1104 33754 34868 33776
rect 1104 33702 9398 33754
rect 9450 33702 9462 33754
rect 9514 33702 9526 33754
rect 9578 33702 9590 33754
rect 9642 33702 9654 33754
rect 9706 33702 17846 33754
rect 17898 33702 17910 33754
rect 17962 33702 17974 33754
rect 18026 33702 18038 33754
rect 18090 33702 18102 33754
rect 18154 33702 26294 33754
rect 26346 33702 26358 33754
rect 26410 33702 26422 33754
rect 26474 33702 26486 33754
rect 26538 33702 26550 33754
rect 26602 33702 34868 33754
rect 1104 33680 34868 33702
rect 10226 33640 10232 33652
rect 10187 33612 10232 33640
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 10318 33504 10324 33516
rect 10279 33476 10324 33504
rect 10318 33464 10324 33476
rect 10376 33464 10382 33516
rect 27614 33504 27620 33516
rect 27575 33476 27620 33504
rect 27614 33464 27620 33476
rect 27672 33464 27678 33516
rect 27798 33436 27804 33448
rect 27759 33408 27804 33436
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 29457 33439 29515 33445
rect 29457 33405 29469 33439
rect 29503 33436 29515 33439
rect 32306 33436 32312 33448
rect 29503 33408 32312 33436
rect 29503 33405 29515 33408
rect 29457 33399 29515 33405
rect 32306 33396 32312 33408
rect 32364 33396 32370 33448
rect 32122 33300 32128 33312
rect 32083 33272 32128 33300
rect 32122 33260 32128 33272
rect 32180 33260 32186 33312
rect 1104 33210 34868 33232
rect 1104 33158 5174 33210
rect 5226 33158 5238 33210
rect 5290 33158 5302 33210
rect 5354 33158 5366 33210
rect 5418 33158 5430 33210
rect 5482 33158 13622 33210
rect 13674 33158 13686 33210
rect 13738 33158 13750 33210
rect 13802 33158 13814 33210
rect 13866 33158 13878 33210
rect 13930 33158 22070 33210
rect 22122 33158 22134 33210
rect 22186 33158 22198 33210
rect 22250 33158 22262 33210
rect 22314 33158 22326 33210
rect 22378 33158 30518 33210
rect 30570 33158 30582 33210
rect 30634 33158 30646 33210
rect 30698 33158 30710 33210
rect 30762 33158 30774 33210
rect 30826 33158 34868 33210
rect 1104 33136 34868 33158
rect 27617 33099 27675 33105
rect 27617 33065 27629 33099
rect 27663 33096 27675 33099
rect 27798 33096 27804 33108
rect 27663 33068 27804 33096
rect 27663 33065 27675 33068
rect 27617 33059 27675 33065
rect 27798 33056 27804 33068
rect 27856 33056 27862 33108
rect 17034 32920 17040 32972
rect 17092 32960 17098 32972
rect 31849 32963 31907 32969
rect 17092 32932 26234 32960
rect 17092 32920 17098 32932
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 18325 32895 18383 32901
rect 18325 32892 18337 32895
rect 18288 32864 18337 32892
rect 18288 32852 18294 32864
rect 18325 32861 18337 32864
rect 18371 32861 18383 32895
rect 26206 32892 26234 32932
rect 31849 32929 31861 32963
rect 31895 32960 31907 32963
rect 32122 32960 32128 32972
rect 31895 32932 32128 32960
rect 31895 32929 31907 32932
rect 31849 32923 31907 32929
rect 32122 32920 32128 32932
rect 32180 32920 32186 32972
rect 27525 32895 27583 32901
rect 27525 32892 27537 32895
rect 26206 32864 27537 32892
rect 18325 32855 18383 32861
rect 27525 32861 27537 32864
rect 27571 32861 27583 32895
rect 27525 32855 27583 32861
rect 29822 32852 29828 32904
rect 29880 32892 29886 32904
rect 30282 32892 30288 32904
rect 29880 32864 30288 32892
rect 29880 32852 29886 32864
rect 30282 32852 30288 32864
rect 30340 32892 30346 32904
rect 31205 32895 31263 32901
rect 31205 32892 31217 32895
rect 30340 32864 31217 32892
rect 30340 32852 30346 32864
rect 31205 32861 31217 32864
rect 31251 32861 31263 32895
rect 31205 32855 31263 32861
rect 31297 32827 31355 32833
rect 31297 32793 31309 32827
rect 31343 32824 31355 32827
rect 32033 32827 32091 32833
rect 32033 32824 32045 32827
rect 31343 32796 32045 32824
rect 31343 32793 31355 32796
rect 31297 32787 31355 32793
rect 32033 32793 32045 32796
rect 32079 32793 32091 32827
rect 33686 32824 33692 32836
rect 33647 32796 33692 32824
rect 32033 32787 32091 32793
rect 33686 32784 33692 32796
rect 33744 32784 33750 32836
rect 1104 32666 34868 32688
rect 1104 32614 9398 32666
rect 9450 32614 9462 32666
rect 9514 32614 9526 32666
rect 9578 32614 9590 32666
rect 9642 32614 9654 32666
rect 9706 32614 17846 32666
rect 17898 32614 17910 32666
rect 17962 32614 17974 32666
rect 18026 32614 18038 32666
rect 18090 32614 18102 32666
rect 18154 32614 26294 32666
rect 26346 32614 26358 32666
rect 26410 32614 26422 32666
rect 26474 32614 26486 32666
rect 26538 32614 26550 32666
rect 26602 32614 34868 32666
rect 1104 32592 34868 32614
rect 20070 32484 20076 32496
rect 20031 32456 20076 32484
rect 20070 32444 20076 32456
rect 20128 32444 20134 32496
rect 18230 32416 18236 32428
rect 18191 32388 18236 32416
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 17954 32308 17960 32360
rect 18012 32348 18018 32360
rect 18417 32351 18475 32357
rect 18417 32348 18429 32351
rect 18012 32320 18429 32348
rect 18012 32308 18018 32320
rect 18417 32317 18429 32320
rect 18463 32317 18475 32351
rect 18417 32311 18475 32317
rect 31573 32351 31631 32357
rect 31573 32317 31585 32351
rect 31619 32348 31631 32351
rect 32125 32351 32183 32357
rect 32125 32348 32137 32351
rect 31619 32320 32137 32348
rect 31619 32317 31631 32320
rect 31573 32311 31631 32317
rect 32125 32317 32137 32320
rect 32171 32317 32183 32351
rect 32306 32348 32312 32360
rect 32267 32320 32312 32348
rect 32125 32311 32183 32317
rect 32306 32308 32312 32320
rect 32364 32308 32370 32360
rect 32585 32351 32643 32357
rect 32585 32317 32597 32351
rect 32631 32317 32643 32351
rect 32585 32311 32643 32317
rect 31846 32240 31852 32292
rect 31904 32280 31910 32292
rect 32600 32280 32628 32311
rect 31904 32252 32628 32280
rect 31904 32240 31910 32252
rect 1104 32122 34868 32144
rect 1104 32070 5174 32122
rect 5226 32070 5238 32122
rect 5290 32070 5302 32122
rect 5354 32070 5366 32122
rect 5418 32070 5430 32122
rect 5482 32070 13622 32122
rect 13674 32070 13686 32122
rect 13738 32070 13750 32122
rect 13802 32070 13814 32122
rect 13866 32070 13878 32122
rect 13930 32070 22070 32122
rect 22122 32070 22134 32122
rect 22186 32070 22198 32122
rect 22250 32070 22262 32122
rect 22314 32070 22326 32122
rect 22378 32070 30518 32122
rect 30570 32070 30582 32122
rect 30634 32070 30646 32122
rect 30698 32070 30710 32122
rect 30762 32070 30774 32122
rect 30826 32070 34868 32122
rect 1104 32048 34868 32070
rect 17954 32008 17960 32020
rect 17915 31980 17960 32008
rect 17954 31968 17960 31980
rect 18012 31968 18018 32020
rect 31665 32011 31723 32017
rect 31665 31977 31677 32011
rect 31711 32008 31723 32011
rect 32306 32008 32312 32020
rect 31711 31980 32312 32008
rect 31711 31977 31723 31980
rect 31665 31971 31723 31977
rect 32306 31968 32312 31980
rect 32364 31968 32370 32020
rect 17034 31832 17040 31884
rect 17092 31872 17098 31884
rect 17586 31872 17592 31884
rect 17092 31844 17592 31872
rect 17092 31832 17098 31844
rect 17586 31832 17592 31844
rect 17644 31832 17650 31884
rect 19518 31832 19524 31884
rect 19576 31872 19582 31884
rect 20717 31875 20775 31881
rect 20717 31872 20729 31875
rect 19576 31844 20729 31872
rect 19576 31832 19582 31844
rect 20717 31841 20729 31844
rect 20763 31841 20775 31875
rect 20717 31835 20775 31841
rect 3418 31764 3424 31816
rect 3476 31804 3482 31816
rect 10962 31804 10968 31816
rect 3476 31776 10968 31804
rect 3476 31764 3482 31776
rect 10962 31764 10968 31776
rect 11020 31764 11026 31816
rect 16298 31764 16304 31816
rect 16356 31804 16362 31816
rect 17865 31807 17923 31813
rect 17865 31804 17877 31807
rect 16356 31776 17877 31804
rect 16356 31764 16362 31776
rect 17865 31773 17877 31776
rect 17911 31773 17923 31807
rect 17865 31767 17923 31773
rect 19613 31807 19671 31813
rect 19613 31773 19625 31807
rect 19659 31804 19671 31807
rect 20073 31807 20131 31813
rect 20073 31804 20085 31807
rect 19659 31776 20085 31804
rect 19659 31773 19671 31776
rect 19613 31767 19671 31773
rect 20073 31773 20085 31776
rect 20119 31773 20131 31807
rect 20073 31767 20131 31773
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31804 26479 31807
rect 26970 31804 26976 31816
rect 26467 31776 26976 31804
rect 26467 31773 26479 31776
rect 26421 31767 26479 31773
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 31573 31807 31631 31813
rect 31573 31773 31585 31807
rect 31619 31804 31631 31807
rect 32030 31804 32036 31816
rect 31619 31776 32036 31804
rect 31619 31773 31631 31776
rect 31573 31767 31631 31773
rect 32030 31764 32036 31776
rect 32088 31764 32094 31816
rect 20254 31736 20260 31748
rect 20215 31708 20260 31736
rect 20254 31696 20260 31708
rect 20312 31696 20318 31748
rect 1104 31578 34868 31600
rect 1104 31526 9398 31578
rect 9450 31526 9462 31578
rect 9514 31526 9526 31578
rect 9578 31526 9590 31578
rect 9642 31526 9654 31578
rect 9706 31526 17846 31578
rect 17898 31526 17910 31578
rect 17962 31526 17974 31578
rect 18026 31526 18038 31578
rect 18090 31526 18102 31578
rect 18154 31526 26294 31578
rect 26346 31526 26358 31578
rect 26410 31526 26422 31578
rect 26474 31526 26486 31578
rect 26538 31526 26550 31578
rect 26602 31526 34868 31578
rect 1104 31504 34868 31526
rect 20254 31464 20260 31476
rect 20215 31436 20260 31464
rect 20254 31424 20260 31436
rect 20312 31424 20318 31476
rect 20162 31328 20168 31340
rect 20123 31300 20168 31328
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 24854 31288 24860 31340
rect 24912 31328 24918 31340
rect 26145 31331 26203 31337
rect 26145 31328 26157 31331
rect 24912 31300 26157 31328
rect 24912 31288 24918 31300
rect 26145 31297 26157 31300
rect 26191 31297 26203 31331
rect 26970 31328 26976 31340
rect 26931 31300 26976 31328
rect 26145 31291 26203 31297
rect 26970 31288 26976 31300
rect 27028 31288 27034 31340
rect 14 31220 20 31272
rect 72 31260 78 31272
rect 10965 31263 11023 31269
rect 72 31232 6914 31260
rect 72 31220 78 31232
rect 6886 31192 6914 31232
rect 10965 31229 10977 31263
rect 11011 31260 11023 31263
rect 11517 31263 11575 31269
rect 11517 31260 11529 31263
rect 11011 31232 11529 31260
rect 11011 31229 11023 31232
rect 10965 31223 11023 31229
rect 11517 31229 11529 31232
rect 11563 31229 11575 31263
rect 11698 31260 11704 31272
rect 11659 31232 11704 31260
rect 11517 31223 11575 31229
rect 11698 31220 11704 31232
rect 11756 31220 11762 31272
rect 11977 31263 12035 31269
rect 11977 31229 11989 31263
rect 12023 31229 12035 31263
rect 11977 31223 12035 31229
rect 26237 31263 26295 31269
rect 26237 31229 26249 31263
rect 26283 31260 26295 31263
rect 27157 31263 27215 31269
rect 27157 31260 27169 31263
rect 26283 31232 27169 31260
rect 26283 31229 26295 31232
rect 26237 31223 26295 31229
rect 27157 31229 27169 31232
rect 27203 31229 27215 31263
rect 27157 31223 27215 31229
rect 27617 31263 27675 31269
rect 27617 31229 27629 31263
rect 27663 31229 27675 31263
rect 27617 31223 27675 31229
rect 11992 31192 12020 31223
rect 6886 31164 12020 31192
rect 26694 31152 26700 31204
rect 26752 31192 26758 31204
rect 27632 31192 27660 31223
rect 26752 31164 27660 31192
rect 26752 31152 26758 31164
rect 1104 31034 34868 31056
rect 1104 30982 5174 31034
rect 5226 30982 5238 31034
rect 5290 30982 5302 31034
rect 5354 30982 5366 31034
rect 5418 30982 5430 31034
rect 5482 30982 13622 31034
rect 13674 30982 13686 31034
rect 13738 30982 13750 31034
rect 13802 30982 13814 31034
rect 13866 30982 13878 31034
rect 13930 30982 22070 31034
rect 22122 30982 22134 31034
rect 22186 30982 22198 31034
rect 22250 30982 22262 31034
rect 22314 30982 22326 31034
rect 22378 30982 30518 31034
rect 30570 30982 30582 31034
rect 30634 30982 30646 31034
rect 30698 30982 30710 31034
rect 30762 30982 30774 31034
rect 30826 30982 34868 31034
rect 1104 30960 34868 30982
rect 11149 30923 11207 30929
rect 11149 30889 11161 30923
rect 11195 30920 11207 30923
rect 11698 30920 11704 30932
rect 11195 30892 11704 30920
rect 11195 30889 11207 30892
rect 11149 30883 11207 30889
rect 11698 30880 11704 30892
rect 11756 30880 11762 30932
rect 2774 30676 2780 30728
rect 2832 30716 2838 30728
rect 2869 30719 2927 30725
rect 2869 30716 2881 30719
rect 2832 30688 2881 30716
rect 2832 30676 2838 30688
rect 2869 30685 2881 30688
rect 2915 30685 2927 30719
rect 2869 30679 2927 30685
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30685 11115 30719
rect 11057 30679 11115 30685
rect 11072 30648 11100 30679
rect 11790 30676 11796 30728
rect 11848 30716 11854 30728
rect 11885 30719 11943 30725
rect 11885 30716 11897 30719
rect 11848 30688 11897 30716
rect 11848 30676 11854 30688
rect 11885 30685 11897 30688
rect 11931 30685 11943 30719
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 11885 30679 11943 30685
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 33962 30716 33968 30728
rect 33923 30688 33968 30716
rect 33962 30676 33968 30688
rect 34020 30676 34026 30728
rect 18230 30648 18236 30660
rect 11072 30620 18236 30648
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 1104 30490 34868 30512
rect 1104 30438 9398 30490
rect 9450 30438 9462 30490
rect 9514 30438 9526 30490
rect 9578 30438 9590 30490
rect 9642 30438 9654 30490
rect 9706 30438 17846 30490
rect 17898 30438 17910 30490
rect 17962 30438 17974 30490
rect 18026 30438 18038 30490
rect 18090 30438 18102 30490
rect 18154 30438 26294 30490
rect 26346 30438 26358 30490
rect 26410 30438 26422 30490
rect 26474 30438 26486 30490
rect 26538 30438 26550 30490
rect 26602 30438 34868 30490
rect 1104 30416 34868 30438
rect 20162 30336 20168 30388
rect 20220 30376 20226 30388
rect 27798 30376 27804 30388
rect 20220 30348 27804 30376
rect 20220 30336 20226 30348
rect 27798 30336 27804 30348
rect 27856 30336 27862 30388
rect 2774 30240 2780 30252
rect 2735 30212 2780 30240
rect 2774 30200 2780 30212
rect 2832 30200 2838 30252
rect 11790 30240 11796 30252
rect 11751 30212 11796 30240
rect 11790 30200 11796 30212
rect 11848 30200 11854 30252
rect 14274 30240 14280 30252
rect 14235 30212 14280 30240
rect 14274 30200 14280 30212
rect 14332 30200 14338 30252
rect 2961 30175 3019 30181
rect 2961 30141 2973 30175
rect 3007 30172 3019 30175
rect 3142 30172 3148 30184
rect 3007 30144 3148 30172
rect 3007 30141 3019 30144
rect 2961 30135 3019 30141
rect 3142 30132 3148 30144
rect 3200 30132 3206 30184
rect 4154 30172 4160 30184
rect 4115 30144 4160 30172
rect 4154 30132 4160 30144
rect 4212 30132 4218 30184
rect 11977 30175 12035 30181
rect 11977 30141 11989 30175
rect 12023 30172 12035 30175
rect 12158 30172 12164 30184
rect 12023 30144 12164 30172
rect 12023 30141 12035 30144
rect 11977 30135 12035 30141
rect 12158 30132 12164 30144
rect 12216 30132 12222 30184
rect 12437 30175 12495 30181
rect 12437 30141 12449 30175
rect 12483 30141 12495 30175
rect 14458 30172 14464 30184
rect 14419 30144 14464 30172
rect 12437 30135 12495 30141
rect 10962 30064 10968 30116
rect 11020 30104 11026 30116
rect 12452 30104 12480 30135
rect 14458 30132 14464 30144
rect 14516 30132 14522 30184
rect 14826 30172 14832 30184
rect 14787 30144 14832 30172
rect 14826 30132 14832 30144
rect 14884 30132 14890 30184
rect 11020 30076 12480 30104
rect 11020 30064 11026 30076
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19429 30039 19487 30045
rect 19429 30036 19441 30039
rect 19392 30008 19441 30036
rect 19392 29996 19398 30008
rect 19429 30005 19441 30008
rect 19475 30005 19487 30039
rect 19429 29999 19487 30005
rect 27062 29996 27068 30048
rect 27120 30036 27126 30048
rect 27157 30039 27215 30045
rect 27157 30036 27169 30039
rect 27120 30008 27169 30036
rect 27120 29996 27126 30008
rect 27157 30005 27169 30008
rect 27203 30005 27215 30039
rect 27157 29999 27215 30005
rect 32306 29996 32312 30048
rect 32364 30036 32370 30048
rect 32953 30039 33011 30045
rect 32953 30036 32965 30039
rect 32364 30008 32965 30036
rect 32364 29996 32370 30008
rect 32953 30005 32965 30008
rect 32999 30005 33011 30039
rect 33778 30036 33784 30048
rect 33739 30008 33784 30036
rect 32953 29999 33011 30005
rect 33778 29996 33784 30008
rect 33836 29996 33842 30048
rect 1104 29946 34868 29968
rect 1104 29894 5174 29946
rect 5226 29894 5238 29946
rect 5290 29894 5302 29946
rect 5354 29894 5366 29946
rect 5418 29894 5430 29946
rect 5482 29894 13622 29946
rect 13674 29894 13686 29946
rect 13738 29894 13750 29946
rect 13802 29894 13814 29946
rect 13866 29894 13878 29946
rect 13930 29894 22070 29946
rect 22122 29894 22134 29946
rect 22186 29894 22198 29946
rect 22250 29894 22262 29946
rect 22314 29894 22326 29946
rect 22378 29894 30518 29946
rect 30570 29894 30582 29946
rect 30634 29894 30646 29946
rect 30698 29894 30710 29946
rect 30762 29894 30774 29946
rect 30826 29894 34868 29946
rect 1104 29872 34868 29894
rect 3142 29832 3148 29844
rect 3103 29804 3148 29832
rect 3142 29792 3148 29804
rect 3200 29792 3206 29844
rect 12158 29832 12164 29844
rect 12119 29804 12164 29832
rect 12158 29792 12164 29804
rect 12216 29792 12222 29844
rect 14458 29832 14464 29844
rect 14419 29804 14464 29832
rect 14458 29792 14464 29804
rect 14516 29792 14522 29844
rect 6886 29736 19840 29764
rect 2958 29588 2964 29640
rect 3016 29628 3022 29640
rect 3237 29631 3295 29637
rect 3237 29628 3249 29631
rect 3016 29600 3249 29628
rect 3016 29588 3022 29600
rect 3237 29597 3249 29600
rect 3283 29597 3295 29631
rect 3237 29591 3295 29597
rect 3418 29520 3424 29572
rect 3476 29560 3482 29572
rect 6886 29560 6914 29736
rect 19334 29696 19340 29708
rect 19295 29668 19340 29696
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 19812 29705 19840 29736
rect 19797 29699 19855 29705
rect 19797 29665 19809 29699
rect 19843 29665 19855 29699
rect 19797 29659 19855 29665
rect 25406 29656 25412 29708
rect 25464 29696 25470 29708
rect 25685 29699 25743 29705
rect 25685 29696 25697 29699
rect 25464 29668 25697 29696
rect 25464 29656 25470 29668
rect 25685 29665 25697 29668
rect 25731 29665 25743 29699
rect 33042 29696 33048 29708
rect 33003 29668 33048 29696
rect 25685 29659 25743 29665
rect 33042 29656 33048 29668
rect 33100 29656 33106 29708
rect 33962 29656 33968 29708
rect 34020 29696 34026 29708
rect 34149 29699 34207 29705
rect 34149 29696 34161 29699
rect 34020 29668 34161 29696
rect 34020 29656 34026 29668
rect 34149 29665 34161 29668
rect 34195 29665 34207 29699
rect 34149 29659 34207 29665
rect 12253 29631 12311 29637
rect 12253 29597 12265 29631
rect 12299 29597 12311 29631
rect 12253 29591 12311 29597
rect 14369 29631 14427 29637
rect 14369 29597 14381 29631
rect 14415 29628 14427 29631
rect 16298 29628 16304 29640
rect 14415 29600 16304 29628
rect 14415 29597 14427 29600
rect 14369 29591 14427 29597
rect 3476 29532 6914 29560
rect 3476 29520 3482 29532
rect 12268 29492 12296 29591
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 25222 29628 25228 29640
rect 25183 29600 25228 29628
rect 25222 29588 25228 29600
rect 25280 29588 25286 29640
rect 27709 29631 27767 29637
rect 27709 29597 27721 29631
rect 27755 29597 27767 29631
rect 27709 29591 27767 29597
rect 28353 29631 28411 29637
rect 28353 29597 28365 29631
rect 28399 29628 28411 29631
rect 29362 29628 29368 29640
rect 28399 29600 29368 29628
rect 28399 29597 28411 29600
rect 28353 29591 28411 29597
rect 19521 29563 19579 29569
rect 19521 29529 19533 29563
rect 19567 29560 19579 29563
rect 19794 29560 19800 29572
rect 19567 29532 19800 29560
rect 19567 29529 19579 29532
rect 19521 29523 19579 29529
rect 19794 29520 19800 29532
rect 19852 29520 19858 29572
rect 25406 29560 25412 29572
rect 25367 29532 25412 29560
rect 25406 29520 25412 29532
rect 25464 29520 25470 29572
rect 27724 29560 27752 29591
rect 29362 29588 29368 29600
rect 29420 29588 29426 29640
rect 33962 29560 33968 29572
rect 26206 29532 27752 29560
rect 33923 29532 33968 29560
rect 19334 29492 19340 29504
rect 12268 29464 19340 29492
rect 19334 29452 19340 29464
rect 19392 29452 19398 29504
rect 20714 29452 20720 29504
rect 20772 29492 20778 29504
rect 26206 29492 26234 29532
rect 33962 29520 33968 29532
rect 34020 29520 34026 29572
rect 20772 29464 26234 29492
rect 20772 29452 20778 29464
rect 27246 29452 27252 29504
rect 27304 29492 27310 29504
rect 27617 29495 27675 29501
rect 27617 29492 27629 29495
rect 27304 29464 27629 29492
rect 27304 29452 27310 29464
rect 27617 29461 27629 29464
rect 27663 29461 27675 29495
rect 27617 29455 27675 29461
rect 1104 29402 34868 29424
rect 1104 29350 9398 29402
rect 9450 29350 9462 29402
rect 9514 29350 9526 29402
rect 9578 29350 9590 29402
rect 9642 29350 9654 29402
rect 9706 29350 17846 29402
rect 17898 29350 17910 29402
rect 17962 29350 17974 29402
rect 18026 29350 18038 29402
rect 18090 29350 18102 29402
rect 18154 29350 26294 29402
rect 26346 29350 26358 29402
rect 26410 29350 26422 29402
rect 26474 29350 26486 29402
rect 26538 29350 26550 29402
rect 26602 29350 34868 29402
rect 1104 29328 34868 29350
rect 2958 29248 2964 29300
rect 3016 29288 3022 29300
rect 18322 29288 18328 29300
rect 3016 29260 18328 29288
rect 3016 29248 3022 29260
rect 18322 29248 18328 29260
rect 18380 29248 18386 29300
rect 19794 29288 19800 29300
rect 19755 29260 19800 29288
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 27246 29220 27252 29232
rect 27207 29192 27252 29220
rect 27246 29180 27252 29192
rect 27304 29180 27310 29232
rect 31205 29223 31263 29229
rect 31205 29189 31217 29223
rect 31251 29220 31263 29223
rect 31662 29220 31668 29232
rect 31251 29192 31668 29220
rect 31251 29189 31263 29192
rect 31205 29183 31263 29189
rect 31662 29180 31668 29192
rect 31720 29180 31726 29232
rect 34146 29220 34152 29232
rect 34107 29192 34152 29220
rect 34146 29180 34152 29192
rect 34204 29180 34210 29232
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 20714 29152 20720 29164
rect 19935 29124 20720 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 25222 29112 25228 29164
rect 25280 29152 25286 29164
rect 26145 29155 26203 29161
rect 26145 29152 26157 29155
rect 25280 29124 26157 29152
rect 25280 29112 25286 29124
rect 26145 29121 26157 29124
rect 26191 29121 26203 29155
rect 27062 29152 27068 29164
rect 27023 29124 27068 29152
rect 26145 29115 26203 29121
rect 27062 29112 27068 29124
rect 27120 29112 27126 29164
rect 29362 29152 29368 29164
rect 29323 29124 29368 29152
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 32306 29152 32312 29164
rect 32267 29124 32312 29152
rect 32306 29112 32312 29124
rect 32364 29112 32370 29164
rect 28442 29084 28448 29096
rect 28403 29056 28448 29084
rect 28442 29044 28448 29056
rect 28500 29044 28506 29096
rect 29546 29084 29552 29096
rect 29507 29056 29552 29084
rect 29546 29044 29552 29056
rect 29604 29044 29610 29096
rect 32490 29084 32496 29096
rect 32451 29056 32496 29084
rect 32490 29044 32496 29056
rect 32548 29044 32554 29096
rect 25498 28948 25504 28960
rect 25459 28920 25504 28948
rect 25498 28908 25504 28920
rect 25556 28908 25562 28960
rect 1104 28858 34868 28880
rect 1104 28806 5174 28858
rect 5226 28806 5238 28858
rect 5290 28806 5302 28858
rect 5354 28806 5366 28858
rect 5418 28806 5430 28858
rect 5482 28806 13622 28858
rect 13674 28806 13686 28858
rect 13738 28806 13750 28858
rect 13802 28806 13814 28858
rect 13866 28806 13878 28858
rect 13930 28806 22070 28858
rect 22122 28806 22134 28858
rect 22186 28806 22198 28858
rect 22250 28806 22262 28858
rect 22314 28806 22326 28858
rect 22378 28806 30518 28858
rect 30570 28806 30582 28858
rect 30634 28806 30646 28858
rect 30698 28806 30710 28858
rect 30762 28806 30774 28858
rect 30826 28806 34868 28858
rect 1104 28784 34868 28806
rect 24949 28747 25007 28753
rect 24949 28713 24961 28747
rect 24995 28744 25007 28747
rect 25406 28744 25412 28756
rect 24995 28716 25412 28744
rect 24995 28713 25007 28716
rect 24949 28707 25007 28713
rect 25406 28704 25412 28716
rect 25464 28704 25470 28756
rect 27893 28747 27951 28753
rect 27893 28713 27905 28747
rect 27939 28744 27951 28747
rect 29546 28744 29552 28756
rect 27939 28716 29552 28744
rect 27939 28713 27951 28716
rect 27893 28707 27951 28713
rect 29546 28704 29552 28716
rect 29604 28704 29610 28756
rect 25498 28608 25504 28620
rect 25459 28580 25504 28608
rect 25498 28568 25504 28580
rect 25556 28568 25562 28620
rect 27341 28611 27399 28617
rect 27341 28577 27353 28611
rect 27387 28608 27399 28611
rect 31570 28608 31576 28620
rect 27387 28580 31576 28608
rect 27387 28577 27399 28580
rect 27341 28571 27399 28577
rect 31570 28568 31576 28580
rect 31628 28568 31634 28620
rect 33502 28608 33508 28620
rect 33463 28580 33508 28608
rect 33502 28568 33508 28580
rect 33560 28568 33566 28620
rect 33778 28568 33784 28620
rect 33836 28608 33842 28620
rect 34149 28611 34207 28617
rect 34149 28608 34161 28611
rect 33836 28580 34161 28608
rect 33836 28568 33842 28580
rect 34149 28577 34161 28580
rect 34195 28577 34207 28611
rect 34149 28571 34207 28577
rect 19702 28500 19708 28552
rect 19760 28540 19766 28552
rect 24854 28540 24860 28552
rect 19760 28512 24860 28540
rect 19760 28500 19766 28512
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 27798 28540 27804 28552
rect 27759 28512 27804 28540
rect 27798 28500 27804 28512
rect 27856 28500 27862 28552
rect 25498 28432 25504 28484
rect 25556 28472 25562 28484
rect 25685 28475 25743 28481
rect 25685 28472 25697 28475
rect 25556 28444 25697 28472
rect 25556 28432 25562 28444
rect 25685 28441 25697 28444
rect 25731 28441 25743 28475
rect 25685 28435 25743 28441
rect 33410 28432 33416 28484
rect 33468 28472 33474 28484
rect 33965 28475 34023 28481
rect 33965 28472 33977 28475
rect 33468 28444 33977 28472
rect 33468 28432 33474 28444
rect 33965 28441 33977 28444
rect 34011 28441 34023 28475
rect 33965 28435 34023 28441
rect 1104 28314 34868 28336
rect 1104 28262 9398 28314
rect 9450 28262 9462 28314
rect 9514 28262 9526 28314
rect 9578 28262 9590 28314
rect 9642 28262 9654 28314
rect 9706 28262 17846 28314
rect 17898 28262 17910 28314
rect 17962 28262 17974 28314
rect 18026 28262 18038 28314
rect 18090 28262 18102 28314
rect 18154 28262 26294 28314
rect 26346 28262 26358 28314
rect 26410 28262 26422 28314
rect 26474 28262 26486 28314
rect 26538 28262 26550 28314
rect 26602 28262 34868 28314
rect 1104 28240 34868 28262
rect 25498 28200 25504 28212
rect 25459 28172 25504 28200
rect 25498 28160 25504 28172
rect 25556 28160 25562 28212
rect 32490 28160 32496 28212
rect 32548 28200 32554 28212
rect 32769 28203 32827 28209
rect 32769 28200 32781 28203
rect 32548 28172 32781 28200
rect 32548 28160 32554 28172
rect 32769 28169 32781 28172
rect 32815 28169 32827 28203
rect 33410 28200 33416 28212
rect 33371 28172 33416 28200
rect 32769 28163 32827 28169
rect 33410 28160 33416 28172
rect 33468 28160 33474 28212
rect 33962 28160 33968 28212
rect 34020 28200 34026 28212
rect 34057 28203 34115 28209
rect 34057 28200 34069 28203
rect 34020 28172 34069 28200
rect 34020 28160 34026 28172
rect 34057 28169 34069 28172
rect 34103 28169 34115 28203
rect 34057 28163 34115 28169
rect 25406 28064 25412 28076
rect 25367 28036 25412 28064
rect 25406 28024 25412 28036
rect 25464 28024 25470 28076
rect 32861 28067 32919 28073
rect 32861 28033 32873 28067
rect 32907 28064 32919 28067
rect 33134 28064 33140 28076
rect 32907 28036 33140 28064
rect 32907 28033 32919 28036
rect 32861 28027 32919 28033
rect 33134 28024 33140 28036
rect 33192 28024 33198 28076
rect 33318 28024 33324 28076
rect 33376 28064 33382 28076
rect 33505 28067 33563 28073
rect 33505 28064 33517 28067
rect 33376 28036 33517 28064
rect 33376 28024 33382 28036
rect 33505 28033 33517 28036
rect 33551 28064 33563 28067
rect 33965 28067 34023 28073
rect 33965 28064 33977 28067
rect 33551 28036 33977 28064
rect 33551 28033 33563 28036
rect 33505 28027 33563 28033
rect 33965 28033 33977 28036
rect 34011 28033 34023 28067
rect 33965 28027 34023 28033
rect 1104 27770 34868 27792
rect 1104 27718 5174 27770
rect 5226 27718 5238 27770
rect 5290 27718 5302 27770
rect 5354 27718 5366 27770
rect 5418 27718 5430 27770
rect 5482 27718 13622 27770
rect 13674 27718 13686 27770
rect 13738 27718 13750 27770
rect 13802 27718 13814 27770
rect 13866 27718 13878 27770
rect 13930 27718 22070 27770
rect 22122 27718 22134 27770
rect 22186 27718 22198 27770
rect 22250 27718 22262 27770
rect 22314 27718 22326 27770
rect 22378 27718 30518 27770
rect 30570 27718 30582 27770
rect 30634 27718 30646 27770
rect 30698 27718 30710 27770
rect 30762 27718 30774 27770
rect 30826 27718 34868 27770
rect 1104 27696 34868 27718
rect 1104 27226 34868 27248
rect 1104 27174 9398 27226
rect 9450 27174 9462 27226
rect 9514 27174 9526 27226
rect 9578 27174 9590 27226
rect 9642 27174 9654 27226
rect 9706 27174 17846 27226
rect 17898 27174 17910 27226
rect 17962 27174 17974 27226
rect 18026 27174 18038 27226
rect 18090 27174 18102 27226
rect 18154 27174 26294 27226
rect 26346 27174 26358 27226
rect 26410 27174 26422 27226
rect 26474 27174 26486 27226
rect 26538 27174 26550 27226
rect 26602 27174 34868 27226
rect 1104 27152 34868 27174
rect 31294 26772 31300 26784
rect 31255 26744 31300 26772
rect 31294 26732 31300 26744
rect 31352 26732 31358 26784
rect 1104 26682 34868 26704
rect 1104 26630 5174 26682
rect 5226 26630 5238 26682
rect 5290 26630 5302 26682
rect 5354 26630 5366 26682
rect 5418 26630 5430 26682
rect 5482 26630 13622 26682
rect 13674 26630 13686 26682
rect 13738 26630 13750 26682
rect 13802 26630 13814 26682
rect 13866 26630 13878 26682
rect 13930 26630 22070 26682
rect 22122 26630 22134 26682
rect 22186 26630 22198 26682
rect 22250 26630 22262 26682
rect 22314 26630 22326 26682
rect 22378 26630 30518 26682
rect 30570 26630 30582 26682
rect 30634 26630 30646 26682
rect 30698 26630 30710 26682
rect 30762 26630 30774 26682
rect 30826 26630 34868 26682
rect 1104 26608 34868 26630
rect 31294 26432 31300 26444
rect 31255 26404 31300 26432
rect 31294 26392 31300 26404
rect 31352 26392 31358 26444
rect 33042 26432 33048 26444
rect 33003 26404 33048 26432
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 8113 26367 8171 26373
rect 8113 26333 8125 26367
rect 8159 26364 8171 26367
rect 8846 26364 8852 26376
rect 8159 26336 8852 26364
rect 8159 26333 8171 26336
rect 8113 26327 8171 26333
rect 8846 26324 8852 26336
rect 8904 26324 8910 26376
rect 29730 26324 29736 26376
rect 29788 26364 29794 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 29788 26336 29837 26364
rect 29788 26324 29794 26336
rect 29825 26333 29837 26336
rect 29871 26333 29883 26367
rect 29825 26327 29883 26333
rect 31481 26299 31539 26305
rect 31481 26265 31493 26299
rect 31527 26296 31539 26299
rect 32214 26296 32220 26308
rect 31527 26268 32220 26296
rect 31527 26265 31539 26268
rect 31481 26259 31539 26265
rect 32214 26256 32220 26268
rect 32272 26256 32278 26308
rect 1104 26138 34868 26160
rect 1104 26086 9398 26138
rect 9450 26086 9462 26138
rect 9514 26086 9526 26138
rect 9578 26086 9590 26138
rect 9642 26086 9654 26138
rect 9706 26086 17846 26138
rect 17898 26086 17910 26138
rect 17962 26086 17974 26138
rect 18026 26086 18038 26138
rect 18090 26086 18102 26138
rect 18154 26086 26294 26138
rect 26346 26086 26358 26138
rect 26410 26086 26422 26138
rect 26474 26086 26486 26138
rect 26538 26086 26550 26138
rect 26602 26086 34868 26138
rect 1104 26064 34868 26086
rect 32214 26024 32220 26036
rect 32175 25996 32220 26024
rect 32214 25984 32220 25996
rect 32272 25984 32278 26036
rect 3602 25916 3608 25968
rect 3660 25956 3666 25968
rect 7837 25959 7895 25965
rect 7837 25956 7849 25959
rect 3660 25928 7849 25956
rect 3660 25916 3666 25928
rect 7837 25925 7849 25928
rect 7883 25925 7895 25959
rect 7837 25919 7895 25925
rect 8846 25916 8852 25968
rect 8904 25956 8910 25968
rect 31573 25959 31631 25965
rect 8904 25928 9720 25956
rect 8904 25916 8910 25928
rect 9692 25897 9720 25928
rect 31573 25925 31585 25959
rect 31619 25956 31631 25959
rect 33042 25956 33048 25968
rect 31619 25928 33048 25956
rect 31619 25925 31631 25928
rect 31573 25919 31631 25925
rect 33042 25916 33048 25928
rect 33100 25916 33106 25968
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 29086 25888 29092 25900
rect 29047 25860 29092 25888
rect 9677 25851 9735 25857
rect 29086 25848 29092 25860
rect 29144 25848 29150 25900
rect 29730 25888 29736 25900
rect 29691 25860 29736 25888
rect 29730 25848 29736 25860
rect 29788 25848 29794 25900
rect 31938 25848 31944 25900
rect 31996 25888 32002 25900
rect 32125 25891 32183 25897
rect 32125 25888 32137 25891
rect 31996 25860 32137 25888
rect 31996 25848 32002 25860
rect 32125 25857 32137 25860
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 9030 25780 9036 25832
rect 9088 25820 9094 25832
rect 9493 25823 9551 25829
rect 9493 25820 9505 25823
rect 9088 25792 9505 25820
rect 9088 25780 9094 25792
rect 9493 25789 9505 25792
rect 9539 25789 9551 25823
rect 9493 25783 9551 25789
rect 29181 25823 29239 25829
rect 29181 25789 29193 25823
rect 29227 25820 29239 25823
rect 29917 25823 29975 25829
rect 29917 25820 29929 25823
rect 29227 25792 29929 25820
rect 29227 25789 29239 25792
rect 29181 25783 29239 25789
rect 29917 25789 29929 25792
rect 29963 25789 29975 25823
rect 29917 25783 29975 25789
rect 9950 25644 9956 25696
rect 10008 25684 10014 25696
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 10008 25656 10149 25684
rect 10008 25644 10014 25656
rect 10137 25653 10149 25656
rect 10183 25653 10195 25687
rect 10137 25647 10195 25653
rect 1104 25594 34868 25616
rect 1104 25542 5174 25594
rect 5226 25542 5238 25594
rect 5290 25542 5302 25594
rect 5354 25542 5366 25594
rect 5418 25542 5430 25594
rect 5482 25542 13622 25594
rect 13674 25542 13686 25594
rect 13738 25542 13750 25594
rect 13802 25542 13814 25594
rect 13866 25542 13878 25594
rect 13930 25542 22070 25594
rect 22122 25542 22134 25594
rect 22186 25542 22198 25594
rect 22250 25542 22262 25594
rect 22314 25542 22326 25594
rect 22378 25542 30518 25594
rect 30570 25542 30582 25594
rect 30634 25542 30646 25594
rect 30698 25542 30710 25594
rect 30762 25542 30774 25594
rect 30826 25542 34868 25594
rect 1104 25520 34868 25542
rect 9030 25480 9036 25492
rect 8991 25452 9036 25480
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 9950 25344 9956 25356
rect 9911 25316 9956 25344
rect 9950 25304 9956 25316
rect 10008 25304 10014 25356
rect 10410 25344 10416 25356
rect 10371 25316 10416 25344
rect 10410 25304 10416 25316
rect 10468 25304 10474 25356
rect 32950 25344 32956 25356
rect 32911 25316 32956 25344
rect 32950 25304 32956 25316
rect 33008 25304 33014 25356
rect 7650 25236 7656 25288
rect 7708 25276 7714 25288
rect 7745 25279 7803 25285
rect 7745 25276 7757 25279
rect 7708 25248 7757 25276
rect 7708 25236 7714 25248
rect 7745 25245 7757 25248
rect 7791 25245 7803 25279
rect 7745 25239 7803 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9306 25276 9312 25288
rect 9171 25248 9312 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9306 25236 9312 25248
rect 9364 25236 9370 25288
rect 31021 25279 31079 25285
rect 31021 25245 31033 25279
rect 31067 25276 31079 25279
rect 31481 25279 31539 25285
rect 31481 25276 31493 25279
rect 31067 25248 31493 25276
rect 31067 25245 31079 25248
rect 31021 25239 31079 25245
rect 31481 25245 31493 25248
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 10134 25208 10140 25220
rect 10095 25180 10140 25208
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 31662 25208 31668 25220
rect 31623 25180 31668 25208
rect 31662 25168 31668 25180
rect 31720 25168 31726 25220
rect 1104 25050 34868 25072
rect 1104 24998 9398 25050
rect 9450 24998 9462 25050
rect 9514 24998 9526 25050
rect 9578 24998 9590 25050
rect 9642 24998 9654 25050
rect 9706 24998 17846 25050
rect 17898 24998 17910 25050
rect 17962 24998 17974 25050
rect 18026 24998 18038 25050
rect 18090 24998 18102 25050
rect 18154 24998 26294 25050
rect 26346 24998 26358 25050
rect 26410 24998 26422 25050
rect 26474 24998 26486 25050
rect 26538 24998 26550 25050
rect 26602 24998 34868 25050
rect 1104 24976 34868 24998
rect 3418 24896 3424 24948
rect 3476 24936 3482 24948
rect 8386 24936 8392 24948
rect 3476 24908 8392 24936
rect 3476 24896 3482 24908
rect 8386 24896 8392 24908
rect 8444 24896 8450 24948
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 10192 24908 10333 24936
rect 10192 24896 10198 24908
rect 10321 24905 10333 24908
rect 10367 24905 10379 24939
rect 10321 24899 10379 24905
rect 31205 24939 31263 24945
rect 31205 24905 31217 24939
rect 31251 24936 31263 24939
rect 31662 24936 31668 24948
rect 31251 24908 31668 24936
rect 31251 24905 31263 24908
rect 31205 24899 31263 24905
rect 31662 24896 31668 24908
rect 31720 24896 31726 24948
rect 7650 24800 7656 24812
rect 7611 24772 7656 24800
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24800 10471 24803
rect 11054 24800 11060 24812
rect 10459 24772 11060 24800
rect 10459 24769 10471 24772
rect 10413 24763 10471 24769
rect 11054 24760 11060 24772
rect 11112 24760 11118 24812
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 25406 24800 25412 24812
rect 18380 24772 25412 24800
rect 18380 24760 18386 24772
rect 25406 24760 25412 24772
rect 25464 24800 25470 24812
rect 27062 24800 27068 24812
rect 25464 24772 27068 24800
rect 25464 24760 25470 24772
rect 27062 24760 27068 24772
rect 27120 24760 27126 24812
rect 31110 24800 31116 24812
rect 31071 24772 31116 24800
rect 31110 24760 31116 24772
rect 31168 24760 31174 24812
rect 7837 24735 7895 24741
rect 7837 24701 7849 24735
rect 7883 24732 7895 24735
rect 8294 24732 8300 24744
rect 7883 24704 8300 24732
rect 7883 24701 7895 24704
rect 7837 24695 7895 24701
rect 8294 24692 8300 24704
rect 8352 24692 8358 24744
rect 8386 24692 8392 24744
rect 8444 24732 8450 24744
rect 8444 24704 8489 24732
rect 8444 24692 8450 24704
rect 32306 24556 32312 24608
rect 32364 24596 32370 24608
rect 32493 24599 32551 24605
rect 32493 24596 32505 24599
rect 32364 24568 32505 24596
rect 32364 24556 32370 24568
rect 32493 24565 32505 24568
rect 32539 24565 32551 24599
rect 32493 24559 32551 24565
rect 1104 24506 34868 24528
rect 1104 24454 5174 24506
rect 5226 24454 5238 24506
rect 5290 24454 5302 24506
rect 5354 24454 5366 24506
rect 5418 24454 5430 24506
rect 5482 24454 13622 24506
rect 13674 24454 13686 24506
rect 13738 24454 13750 24506
rect 13802 24454 13814 24506
rect 13866 24454 13878 24506
rect 13930 24454 22070 24506
rect 22122 24454 22134 24506
rect 22186 24454 22198 24506
rect 22250 24454 22262 24506
rect 22314 24454 22326 24506
rect 22378 24454 30518 24506
rect 30570 24454 30582 24506
rect 30634 24454 30646 24506
rect 30698 24454 30710 24506
rect 30762 24454 30774 24506
rect 30826 24454 34868 24506
rect 1104 24432 34868 24454
rect 8294 24392 8300 24404
rect 8255 24364 8300 24392
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24188 8447 24191
rect 11054 24188 11060 24200
rect 8435 24160 11060 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 29822 24188 29828 24200
rect 26206 24160 29828 24188
rect 19610 24080 19616 24132
rect 19668 24120 19674 24132
rect 19705 24123 19763 24129
rect 19705 24120 19717 24123
rect 19668 24092 19717 24120
rect 19668 24080 19674 24092
rect 19705 24089 19717 24092
rect 19751 24089 19763 24123
rect 19705 24083 19763 24089
rect 19981 24055 20039 24061
rect 19981 24021 19993 24055
rect 20027 24052 20039 24055
rect 26206 24052 26234 24160
rect 29822 24148 29828 24160
rect 29880 24148 29886 24200
rect 30837 24191 30895 24197
rect 30837 24157 30849 24191
rect 30883 24188 30895 24191
rect 30926 24188 30932 24200
rect 30883 24160 30932 24188
rect 30883 24157 30895 24160
rect 30837 24151 30895 24157
rect 30926 24148 30932 24160
rect 30984 24148 30990 24200
rect 32030 24148 32036 24200
rect 32088 24188 32094 24200
rect 32125 24191 32183 24197
rect 32125 24188 32137 24191
rect 32088 24160 32137 24188
rect 32088 24148 32094 24160
rect 32125 24157 32137 24160
rect 32171 24157 32183 24191
rect 32766 24188 32772 24200
rect 32727 24160 32772 24188
rect 32125 24151 32183 24157
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 29914 24052 29920 24064
rect 20027 24024 26234 24052
rect 29875 24024 29920 24052
rect 20027 24021 20039 24024
rect 19981 24015 20039 24021
rect 29914 24012 29920 24024
rect 29972 24012 29978 24064
rect 32217 24055 32275 24061
rect 32217 24021 32229 24055
rect 32263 24052 32275 24055
rect 32490 24052 32496 24064
rect 32263 24024 32496 24052
rect 32263 24021 32275 24024
rect 32217 24015 32275 24021
rect 32490 24012 32496 24024
rect 32548 24012 32554 24064
rect 1104 23962 34868 23984
rect 1104 23910 9398 23962
rect 9450 23910 9462 23962
rect 9514 23910 9526 23962
rect 9578 23910 9590 23962
rect 9642 23910 9654 23962
rect 9706 23910 17846 23962
rect 17898 23910 17910 23962
rect 17962 23910 17974 23962
rect 18026 23910 18038 23962
rect 18090 23910 18102 23962
rect 18154 23910 26294 23962
rect 26346 23910 26358 23962
rect 26410 23910 26422 23962
rect 26474 23910 26486 23962
rect 26538 23910 26550 23962
rect 26602 23910 34868 23962
rect 1104 23888 34868 23910
rect 17497 23851 17555 23857
rect 17497 23817 17509 23851
rect 17543 23817 17555 23851
rect 17497 23811 17555 23817
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 16574 23712 16580 23724
rect 2004 23684 16580 23712
rect 2004 23672 2010 23684
rect 16574 23672 16580 23684
rect 16632 23712 16638 23724
rect 17313 23715 17371 23721
rect 17313 23712 17325 23715
rect 16632 23684 17325 23712
rect 16632 23672 16638 23684
rect 17313 23681 17325 23684
rect 17359 23681 17371 23715
rect 17512 23712 17540 23811
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23780 18291 23783
rect 18322 23780 18328 23792
rect 18279 23752 18328 23780
rect 18279 23749 18291 23752
rect 18233 23743 18291 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 29914 23780 29920 23792
rect 29875 23752 29920 23780
rect 29914 23740 29920 23752
rect 29972 23740 29978 23792
rect 32490 23780 32496 23792
rect 32451 23752 32496 23780
rect 32490 23740 32496 23752
rect 32548 23740 32554 23792
rect 34146 23780 34152 23792
rect 34107 23752 34152 23780
rect 34146 23740 34152 23752
rect 34204 23740 34210 23792
rect 17957 23715 18015 23721
rect 17957 23712 17969 23715
rect 17512 23684 17969 23712
rect 17313 23675 17371 23681
rect 17957 23681 17969 23684
rect 18003 23712 18015 23715
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 18003 23684 19257 23712
rect 18003 23681 18015 23684
rect 17957 23675 18015 23681
rect 19245 23681 19257 23684
rect 19291 23712 19303 23715
rect 19610 23712 19616 23724
rect 19291 23684 19616 23712
rect 19291 23681 19303 23684
rect 19245 23675 19303 23681
rect 19610 23672 19616 23684
rect 19668 23712 19674 23724
rect 19978 23712 19984 23724
rect 19668 23684 19984 23712
rect 19668 23672 19674 23684
rect 19978 23672 19984 23684
rect 20036 23712 20042 23724
rect 20165 23715 20223 23721
rect 20165 23712 20177 23715
rect 20036 23684 20177 23712
rect 20036 23672 20042 23684
rect 20165 23681 20177 23684
rect 20211 23681 20223 23715
rect 32306 23712 32312 23724
rect 32267 23684 32312 23712
rect 20165 23675 20223 23681
rect 32306 23672 32312 23684
rect 32364 23672 32370 23724
rect 29730 23644 29736 23656
rect 29691 23616 29736 23644
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 30193 23647 30251 23653
rect 30193 23613 30205 23647
rect 30239 23613 30251 23647
rect 30193 23607 30251 23613
rect 19352 23548 26234 23576
rect 19352 23520 19380 23548
rect 19334 23508 19340 23520
rect 19295 23480 19340 23508
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 20441 23511 20499 23517
rect 20441 23477 20453 23511
rect 20487 23508 20499 23511
rect 20714 23508 20720 23520
rect 20487 23480 20720 23508
rect 20487 23477 20499 23480
rect 20441 23471 20499 23477
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 26206 23508 26234 23548
rect 29178 23536 29184 23588
rect 29236 23576 29242 23588
rect 30208 23576 30236 23607
rect 29236 23548 30236 23576
rect 29236 23536 29242 23548
rect 32030 23508 32036 23520
rect 26206 23480 32036 23508
rect 32030 23468 32036 23480
rect 32088 23468 32094 23520
rect 1104 23418 34868 23440
rect 1104 23366 5174 23418
rect 5226 23366 5238 23418
rect 5290 23366 5302 23418
rect 5354 23366 5366 23418
rect 5418 23366 5430 23418
rect 5482 23366 13622 23418
rect 13674 23366 13686 23418
rect 13738 23366 13750 23418
rect 13802 23366 13814 23418
rect 13866 23366 13878 23418
rect 13930 23366 22070 23418
rect 22122 23366 22134 23418
rect 22186 23366 22198 23418
rect 22250 23366 22262 23418
rect 22314 23366 22326 23418
rect 22378 23366 30518 23418
rect 30570 23366 30582 23418
rect 30634 23366 30646 23418
rect 30698 23366 30710 23418
rect 30762 23366 30774 23418
rect 30826 23366 34868 23418
rect 1104 23344 34868 23366
rect 29730 23264 29736 23316
rect 29788 23304 29794 23316
rect 29825 23307 29883 23313
rect 29825 23304 29837 23307
rect 29788 23276 29837 23304
rect 29788 23264 29794 23276
rect 29825 23273 29837 23276
rect 29871 23273 29883 23307
rect 29825 23267 29883 23273
rect 30926 23236 30932 23248
rect 30852 23208 30932 23236
rect 30852 23177 30880 23208
rect 30926 23196 30932 23208
rect 30984 23196 30990 23248
rect 30837 23171 30895 23177
rect 30837 23137 30849 23171
rect 30883 23137 30895 23171
rect 32674 23168 32680 23180
rect 32635 23140 32680 23168
rect 30837 23131 30895 23137
rect 32674 23128 32680 23140
rect 32732 23128 32738 23180
rect 19978 23100 19984 23112
rect 19939 23072 19984 23100
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 33134 23100 33140 23112
rect 33095 23072 33140 23100
rect 33134 23060 33140 23072
rect 33192 23060 33198 23112
rect 30834 22992 30840 23044
rect 30892 23032 30898 23044
rect 31021 23035 31079 23041
rect 31021 23032 31033 23035
rect 30892 23004 31033 23032
rect 30892 22992 30898 23004
rect 31021 23001 31033 23004
rect 31067 23001 31079 23035
rect 31021 22995 31079 23001
rect 19702 22964 19708 22976
rect 19663 22936 19708 22964
rect 19702 22924 19708 22936
rect 19760 22924 19766 22976
rect 32490 22924 32496 22976
rect 32548 22964 32554 22976
rect 33229 22967 33287 22973
rect 33229 22964 33241 22967
rect 32548 22936 33241 22964
rect 32548 22924 32554 22936
rect 33229 22933 33241 22936
rect 33275 22933 33287 22967
rect 33229 22927 33287 22933
rect 1104 22874 34868 22896
rect 1104 22822 9398 22874
rect 9450 22822 9462 22874
rect 9514 22822 9526 22874
rect 9578 22822 9590 22874
rect 9642 22822 9654 22874
rect 9706 22822 17846 22874
rect 17898 22822 17910 22874
rect 17962 22822 17974 22874
rect 18026 22822 18038 22874
rect 18090 22822 18102 22874
rect 18154 22822 26294 22874
rect 26346 22822 26358 22874
rect 26410 22822 26422 22874
rect 26474 22822 26486 22874
rect 26538 22822 26550 22874
rect 26602 22822 34868 22874
rect 1104 22800 34868 22822
rect 30834 22760 30840 22772
rect 30795 22732 30840 22760
rect 30834 22720 30840 22732
rect 30892 22720 30898 22772
rect 32490 22692 32496 22704
rect 32451 22664 32496 22692
rect 32490 22652 32496 22664
rect 32548 22652 32554 22704
rect 34146 22692 34152 22704
rect 34107 22664 34152 22692
rect 34146 22652 34152 22664
rect 34204 22652 34210 22704
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 30745 22627 30803 22633
rect 30745 22624 30757 22627
rect 30432 22596 30757 22624
rect 30432 22584 30438 22596
rect 30745 22593 30757 22596
rect 30791 22624 30803 22627
rect 31110 22624 31116 22636
rect 30791 22596 31116 22624
rect 30791 22593 30803 22596
rect 30745 22587 30803 22593
rect 31110 22584 31116 22596
rect 31168 22584 31174 22636
rect 32309 22559 32367 22565
rect 32309 22525 32321 22559
rect 32355 22556 32367 22559
rect 32766 22556 32772 22568
rect 32355 22528 32772 22556
rect 32355 22525 32367 22528
rect 32309 22519 32367 22525
rect 32766 22516 32772 22528
rect 32824 22516 32830 22568
rect 1104 22330 34868 22352
rect 1104 22278 5174 22330
rect 5226 22278 5238 22330
rect 5290 22278 5302 22330
rect 5354 22278 5366 22330
rect 5418 22278 5430 22330
rect 5482 22278 13622 22330
rect 13674 22278 13686 22330
rect 13738 22278 13750 22330
rect 13802 22278 13814 22330
rect 13866 22278 13878 22330
rect 13930 22278 22070 22330
rect 22122 22278 22134 22330
rect 22186 22278 22198 22330
rect 22250 22278 22262 22330
rect 22314 22278 22326 22330
rect 22378 22278 30518 22330
rect 30570 22278 30582 22330
rect 30634 22278 30646 22330
rect 30698 22278 30710 22330
rect 30762 22278 30774 22330
rect 30826 22278 34868 22330
rect 1104 22256 34868 22278
rect 1104 21786 34868 21808
rect 1104 21734 9398 21786
rect 9450 21734 9462 21786
rect 9514 21734 9526 21786
rect 9578 21734 9590 21786
rect 9642 21734 9654 21786
rect 9706 21734 17846 21786
rect 17898 21734 17910 21786
rect 17962 21734 17974 21786
rect 18026 21734 18038 21786
rect 18090 21734 18102 21786
rect 18154 21734 26294 21786
rect 26346 21734 26358 21786
rect 26410 21734 26422 21786
rect 26474 21734 26486 21786
rect 26538 21734 26550 21786
rect 26602 21734 34868 21786
rect 1104 21712 34868 21734
rect 17678 21536 17684 21548
rect 17639 21508 17684 21536
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 17000 21440 17509 21468
rect 17000 21428 17006 21440
rect 17497 21437 17509 21440
rect 17543 21468 17555 21471
rect 23474 21468 23480 21480
rect 17543 21440 23480 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 1104 21242 34868 21264
rect 1104 21190 5174 21242
rect 5226 21190 5238 21242
rect 5290 21190 5302 21242
rect 5354 21190 5366 21242
rect 5418 21190 5430 21242
rect 5482 21190 13622 21242
rect 13674 21190 13686 21242
rect 13738 21190 13750 21242
rect 13802 21190 13814 21242
rect 13866 21190 13878 21242
rect 13930 21190 22070 21242
rect 22122 21190 22134 21242
rect 22186 21190 22198 21242
rect 22250 21190 22262 21242
rect 22314 21190 22326 21242
rect 22378 21190 30518 21242
rect 30570 21190 30582 21242
rect 30634 21190 30646 21242
rect 30698 21190 30710 21242
rect 30762 21190 30774 21242
rect 30826 21190 34868 21242
rect 1104 21168 34868 21190
rect 17218 20884 17224 20936
rect 17276 20924 17282 20936
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 17276 20896 17325 20924
rect 17276 20884 17282 20896
rect 17313 20893 17325 20896
rect 17359 20924 17371 20927
rect 17678 20924 17684 20936
rect 17359 20896 17684 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17678 20884 17684 20896
rect 17736 20884 17742 20936
rect 28350 20924 28356 20936
rect 28311 20896 28356 20924
rect 28350 20884 28356 20896
rect 28408 20884 28414 20936
rect 29546 20924 29552 20936
rect 29507 20896 29552 20924
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 17586 20788 17592 20800
rect 17547 20760 17592 20788
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 1104 20698 34868 20720
rect 1104 20646 9398 20698
rect 9450 20646 9462 20698
rect 9514 20646 9526 20698
rect 9578 20646 9590 20698
rect 9642 20646 9654 20698
rect 9706 20646 17846 20698
rect 17898 20646 17910 20698
rect 17962 20646 17974 20698
rect 18026 20646 18038 20698
rect 18090 20646 18102 20698
rect 18154 20646 26294 20698
rect 26346 20646 26358 20698
rect 26410 20646 26422 20698
rect 26474 20646 26486 20698
rect 26538 20646 26550 20698
rect 26602 20646 34868 20698
rect 1104 20624 34868 20646
rect 10318 20516 10324 20528
rect 9232 20488 10324 20516
rect 9232 20457 9260 20488
rect 10318 20476 10324 20488
rect 10376 20516 10382 20528
rect 30193 20519 30251 20525
rect 10376 20488 18552 20516
rect 10376 20476 10382 20488
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16574 20448 16580 20460
rect 15979 20420 16580 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16574 20408 16580 20420
rect 16632 20448 16638 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16632 20420 16957 20448
rect 16632 20408 16638 20420
rect 16945 20417 16957 20420
rect 16991 20448 17003 20451
rect 17034 20448 17040 20460
rect 16991 20420 17040 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 18524 20389 18552 20488
rect 30193 20485 30205 20519
rect 30239 20516 30251 20519
rect 32950 20516 32956 20528
rect 30239 20488 32956 20516
rect 30239 20485 30251 20488
rect 30193 20479 30251 20485
rect 32950 20476 32956 20488
rect 33008 20476 33014 20528
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 27709 20451 27767 20457
rect 27709 20448 27721 20451
rect 20772 20420 27721 20448
rect 20772 20408 20778 20420
rect 27709 20417 27721 20420
rect 27755 20417 27767 20451
rect 28350 20448 28356 20460
rect 28311 20420 28356 20448
rect 27709 20411 27767 20417
rect 28350 20408 28356 20420
rect 28408 20408 28414 20460
rect 18509 20383 18567 20389
rect 18509 20349 18521 20383
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 27801 20383 27859 20389
rect 27801 20349 27813 20383
rect 27847 20380 27859 20383
rect 28537 20383 28595 20389
rect 28537 20380 28549 20383
rect 27847 20352 28549 20380
rect 27847 20349 27859 20352
rect 27801 20343 27859 20349
rect 28537 20349 28549 20352
rect 28583 20349 28595 20383
rect 28537 20343 28595 20349
rect 18524 20312 18552 20343
rect 29086 20312 29092 20324
rect 18524 20284 29092 20312
rect 29086 20272 29092 20284
rect 29144 20272 29150 20324
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8536 20216 8585 20244
rect 8536 20204 8542 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8720 20216 9137 20244
rect 8720 20204 8726 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 16117 20247 16175 20253
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16850 20244 16856 20256
rect 16163 20216 16856 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 24578 20204 24584 20256
rect 24636 20244 24642 20256
rect 24673 20247 24731 20253
rect 24673 20244 24685 20247
rect 24636 20216 24685 20244
rect 24636 20204 24642 20216
rect 24673 20213 24685 20216
rect 24719 20213 24731 20247
rect 24673 20207 24731 20213
rect 1104 20154 34868 20176
rect 1104 20102 5174 20154
rect 5226 20102 5238 20154
rect 5290 20102 5302 20154
rect 5354 20102 5366 20154
rect 5418 20102 5430 20154
rect 5482 20102 13622 20154
rect 13674 20102 13686 20154
rect 13738 20102 13750 20154
rect 13802 20102 13814 20154
rect 13866 20102 13878 20154
rect 13930 20102 22070 20154
rect 22122 20102 22134 20154
rect 22186 20102 22198 20154
rect 22250 20102 22262 20154
rect 22314 20102 22326 20154
rect 22378 20102 30518 20154
rect 30570 20102 30582 20154
rect 30634 20102 30646 20154
rect 30698 20102 30710 20154
rect 30762 20102 30774 20154
rect 30826 20102 34868 20154
rect 1104 20080 34868 20102
rect 16298 20040 16304 20052
rect 16259 20012 16304 20040
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 17586 19932 17592 19984
rect 17644 19972 17650 19984
rect 17644 19944 26234 19972
rect 17644 19932 17650 19944
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 6886 19876 11529 19904
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 6886 19768 6914 19876
rect 11517 19873 11529 19876
rect 11563 19873 11575 19907
rect 17034 19904 17040 19916
rect 16995 19876 17040 19904
rect 11517 19867 11575 19873
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 24578 19904 24584 19916
rect 24539 19876 24584 19904
rect 24578 19864 24584 19876
rect 24636 19864 24642 19916
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 9180 19808 9413 19836
rect 9180 19796 9186 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 10643 19808 11069 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 11057 19805 11069 19808
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 17402 19836 17408 19848
rect 17359 19808 17408 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 26206 19836 26234 19944
rect 29546 19904 29552 19916
rect 29507 19876 29552 19904
rect 29546 19864 29552 19876
rect 29604 19864 29610 19916
rect 28813 19839 28871 19845
rect 28813 19836 28825 19839
rect 26206 19808 28825 19836
rect 28813 19805 28825 19808
rect 28859 19805 28871 19839
rect 28813 19799 28871 19805
rect 3568 19740 6914 19768
rect 11241 19771 11299 19777
rect 3568 19728 3574 19740
rect 11241 19737 11253 19771
rect 11287 19768 11299 19771
rect 11606 19768 11612 19780
rect 11287 19740 11612 19768
rect 11287 19737 11299 19740
rect 11241 19731 11299 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 16209 19771 16267 19777
rect 16209 19737 16221 19771
rect 16255 19768 16267 19771
rect 16850 19768 16856 19780
rect 16255 19740 16856 19768
rect 16255 19737 16267 19740
rect 16209 19731 16267 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 24302 19728 24308 19780
rect 24360 19768 24366 19780
rect 24765 19771 24823 19777
rect 24765 19768 24777 19771
rect 24360 19740 24777 19768
rect 24360 19728 24366 19740
rect 24765 19737 24777 19740
rect 24811 19737 24823 19771
rect 24765 19731 24823 19737
rect 26421 19771 26479 19777
rect 26421 19737 26433 19771
rect 26467 19737 26479 19771
rect 26421 19731 26479 19737
rect 28905 19771 28963 19777
rect 28905 19737 28917 19771
rect 28951 19768 28963 19771
rect 29733 19771 29791 19777
rect 29733 19768 29745 19771
rect 28951 19740 29745 19768
rect 28951 19737 28963 19740
rect 28905 19731 28963 19737
rect 29733 19737 29745 19740
rect 29779 19737 29791 19771
rect 31386 19768 31392 19780
rect 31347 19740 31392 19768
rect 29733 19731 29791 19737
rect 26436 19700 26464 19731
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 31754 19700 31760 19712
rect 26436 19672 31760 19700
rect 31754 19660 31760 19672
rect 31812 19660 31818 19712
rect 1104 19610 34868 19632
rect 1104 19558 9398 19610
rect 9450 19558 9462 19610
rect 9514 19558 9526 19610
rect 9578 19558 9590 19610
rect 9642 19558 9654 19610
rect 9706 19558 17846 19610
rect 17898 19558 17910 19610
rect 17962 19558 17974 19610
rect 18026 19558 18038 19610
rect 18090 19558 18102 19610
rect 18154 19558 26294 19610
rect 26346 19558 26358 19610
rect 26410 19558 26422 19610
rect 26474 19558 26486 19610
rect 26538 19558 26550 19610
rect 26602 19558 34868 19610
rect 1104 19536 34868 19558
rect 11606 19496 11612 19508
rect 11567 19468 11612 19496
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 20162 19496 20168 19508
rect 17972 19468 20168 19496
rect 8662 19428 8668 19440
rect 8623 19400 8668 19428
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 17126 19428 17132 19440
rect 16546 19400 17132 19428
rect 8478 19360 8484 19372
rect 8439 19332 8484 19360
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 10318 19360 10324 19372
rect 10279 19332 10324 19360
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 16546 19360 16574 19400
rect 17126 19388 17132 19400
rect 17184 19388 17190 19440
rect 17972 19428 18000 19468
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 24302 19496 24308 19508
rect 24263 19468 24308 19496
rect 24302 19456 24308 19468
rect 24360 19456 24366 19508
rect 17236 19400 18000 19428
rect 18049 19431 18107 19437
rect 16850 19360 16856 19372
rect 11747 19332 16574 19360
rect 16763 19332 16856 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 16868 19224 16896 19320
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 17092 19264 17141 19292
rect 17092 19252 17098 19264
rect 17129 19261 17141 19264
rect 17175 19292 17187 19295
rect 17236 19292 17264 19400
rect 18049 19397 18061 19431
rect 18095 19428 18107 19431
rect 18230 19428 18236 19440
rect 18095 19400 18236 19428
rect 18095 19397 18107 19400
rect 18049 19391 18107 19397
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 18874 19388 18880 19440
rect 18932 19428 18938 19440
rect 18969 19431 19027 19437
rect 18969 19428 18981 19431
rect 18932 19400 18981 19428
rect 18932 19388 18938 19400
rect 18969 19397 18981 19400
rect 19015 19428 19027 19431
rect 30374 19428 30380 19440
rect 19015 19400 30380 19428
rect 19015 19397 19027 19400
rect 18969 19391 19027 19397
rect 30374 19388 30380 19400
rect 30432 19388 30438 19440
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17460 19332 17785 19360
rect 17460 19320 17466 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 18690 19360 18696 19372
rect 17773 19323 17831 19329
rect 17880 19332 18696 19360
rect 17175 19264 17264 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17494 19224 17500 19236
rect 16868 19196 17500 19224
rect 17494 19184 17500 19196
rect 17552 19224 17558 19236
rect 17880 19224 17908 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 23474 19320 23480 19372
rect 23532 19360 23538 19372
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23532 19332 24225 19360
rect 23532 19320 23538 19332
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 33042 19292 33048 19304
rect 33003 19264 33048 19292
rect 33042 19252 33048 19264
rect 33100 19252 33106 19304
rect 33226 19252 33232 19304
rect 33284 19292 33290 19304
rect 33965 19295 34023 19301
rect 33965 19292 33977 19295
rect 33284 19264 33977 19292
rect 33284 19252 33290 19264
rect 33965 19261 33977 19264
rect 34011 19261 34023 19295
rect 34146 19292 34152 19304
rect 34107 19264 34152 19292
rect 33965 19255 34023 19261
rect 34146 19252 34152 19264
rect 34204 19252 34210 19304
rect 17552 19196 17908 19224
rect 17552 19184 17558 19196
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 6365 19159 6423 19165
rect 6365 19156 6377 19159
rect 6328 19128 6377 19156
rect 6328 19116 6334 19128
rect 6365 19125 6377 19128
rect 6411 19125 6423 19159
rect 6365 19119 6423 19125
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10284 19128 10793 19156
rect 10284 19116 10290 19128
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 10781 19119 10839 19125
rect 1104 19066 34868 19088
rect 1104 19014 5174 19066
rect 5226 19014 5238 19066
rect 5290 19014 5302 19066
rect 5354 19014 5366 19066
rect 5418 19014 5430 19066
rect 5482 19014 13622 19066
rect 13674 19014 13686 19066
rect 13738 19014 13750 19066
rect 13802 19014 13814 19066
rect 13866 19014 13878 19066
rect 13930 19014 22070 19066
rect 22122 19014 22134 19066
rect 22186 19014 22198 19066
rect 22250 19014 22262 19066
rect 22314 19014 22326 19066
rect 22378 19014 30518 19066
rect 30570 19014 30582 19066
rect 30634 19014 30646 19066
rect 30698 19014 30710 19066
rect 30762 19014 30774 19066
rect 30826 19014 34868 19066
rect 1104 18992 34868 19014
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 9364 18924 17264 18952
rect 9364 18912 9370 18924
rect 17236 18884 17264 18924
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 17368 18924 17509 18952
rect 17368 18912 17374 18924
rect 17497 18921 17509 18924
rect 17543 18952 17555 18955
rect 17678 18952 17684 18964
rect 17543 18924 17684 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 33226 18952 33232 18964
rect 33187 18924 33232 18952
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 33965 18955 34023 18961
rect 33965 18921 33977 18955
rect 34011 18952 34023 18955
rect 34146 18952 34152 18964
rect 34011 18924 34152 18952
rect 34011 18921 34023 18924
rect 33965 18915 34023 18921
rect 34146 18912 34152 18924
rect 34204 18912 34210 18964
rect 19150 18884 19156 18896
rect 9140 18856 16574 18884
rect 17236 18856 19156 18884
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 9140 18757 9168 18856
rect 10226 18816 10232 18828
rect 10187 18788 10232 18816
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 10686 18816 10692 18828
rect 10647 18788 10692 18816
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 16546 18816 16574 18856
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 31662 18884 31668 18896
rect 29012 18856 31668 18884
rect 19334 18816 19340 18828
rect 16546 18788 19340 18816
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 29012 18825 29040 18856
rect 31662 18844 31668 18856
rect 31720 18844 31726 18896
rect 28997 18819 29055 18825
rect 28997 18785 29009 18819
rect 29043 18785 29055 18819
rect 28997 18779 29055 18785
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 5132 18720 5273 18748
rect 5132 18708 5138 18720
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9364 18720 9597 18748
rect 9364 18708 9370 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 17218 18748 17224 18760
rect 16807 18720 17224 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 27154 18748 27160 18760
rect 27115 18720 27160 18748
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18748 31723 18751
rect 32030 18748 32036 18760
rect 31711 18720 32036 18748
rect 31711 18717 31723 18720
rect 31665 18711 31723 18717
rect 32030 18708 32036 18720
rect 32088 18708 32094 18760
rect 32122 18708 32128 18760
rect 32180 18748 32186 18760
rect 32309 18751 32367 18757
rect 32309 18748 32321 18751
rect 32180 18720 32321 18748
rect 32180 18708 32186 18720
rect 32309 18717 32321 18720
rect 32355 18717 32367 18751
rect 32309 18711 32367 18717
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18748 33195 18751
rect 33318 18748 33324 18760
rect 33183 18720 33324 18748
rect 33183 18717 33195 18720
rect 33137 18711 33195 18717
rect 6457 18683 6515 18689
rect 6457 18649 6469 18683
rect 6503 18680 6515 18683
rect 6638 18680 6644 18692
rect 6503 18652 6644 18680
rect 6503 18649 6515 18652
rect 6457 18643 6515 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 8110 18680 8116 18692
rect 8071 18652 8116 18680
rect 8110 18640 8116 18652
rect 8168 18640 8174 18692
rect 9677 18683 9735 18689
rect 8956 18652 9444 18680
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 8956 18612 8984 18652
rect 3476 18584 8984 18612
rect 3476 18572 3482 18584
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9416 18612 9444 18652
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 10413 18683 10471 18689
rect 10413 18680 10425 18683
rect 9723 18652 10425 18680
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 10413 18649 10425 18652
rect 10459 18649 10471 18683
rect 17402 18680 17408 18692
rect 17363 18652 17408 18680
rect 10413 18643 10471 18649
rect 17402 18640 17408 18652
rect 17460 18680 17466 18692
rect 18325 18683 18383 18689
rect 18325 18680 18337 18683
rect 17460 18652 18337 18680
rect 17460 18640 17466 18652
rect 18325 18649 18337 18652
rect 18371 18649 18383 18683
rect 27338 18680 27344 18692
rect 27299 18652 27344 18680
rect 18325 18643 18383 18649
rect 27338 18640 27344 18652
rect 27396 18640 27402 18692
rect 33152 18680 33180 18711
rect 33318 18708 33324 18720
rect 33376 18748 33382 18760
rect 33778 18748 33784 18760
rect 33376 18720 33784 18748
rect 33376 18708 33382 18720
rect 33778 18708 33784 18720
rect 33836 18708 33842 18760
rect 31588 18652 33180 18680
rect 10686 18612 10692 18624
rect 9088 18584 9133 18612
rect 9416 18584 10692 18612
rect 9088 18572 9094 18584
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 16482 18612 16488 18624
rect 11112 18584 16488 18612
rect 11112 18572 11118 18584
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 17828 18584 18613 18612
rect 17828 18572 17834 18584
rect 18601 18581 18613 18584
rect 18647 18612 18659 18615
rect 31588 18612 31616 18652
rect 18647 18584 31616 18612
rect 31757 18615 31815 18621
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 31757 18581 31769 18615
rect 31803 18612 31815 18615
rect 32306 18612 32312 18624
rect 31803 18584 32312 18612
rect 31803 18581 31815 18584
rect 31757 18575 31815 18581
rect 32306 18572 32312 18584
rect 32364 18572 32370 18624
rect 1104 18522 34868 18544
rect 1104 18470 9398 18522
rect 9450 18470 9462 18522
rect 9514 18470 9526 18522
rect 9578 18470 9590 18522
rect 9642 18470 9654 18522
rect 9706 18470 17846 18522
rect 17898 18470 17910 18522
rect 17962 18470 17974 18522
rect 18026 18470 18038 18522
rect 18090 18470 18102 18522
rect 18154 18470 26294 18522
rect 26346 18470 26358 18522
rect 26410 18470 26422 18522
rect 26474 18470 26486 18522
rect 26538 18470 26550 18522
rect 26602 18470 34868 18522
rect 1104 18448 34868 18470
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 16942 18408 16948 18420
rect 6788 18380 16948 18408
rect 6788 18368 6794 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 6748 18281 6776 18368
rect 10965 18343 11023 18349
rect 10965 18340 10977 18343
rect 6886 18312 10977 18340
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18241 6791 18275
rect 6733 18235 6791 18241
rect 3418 18164 3424 18216
rect 3476 18204 3482 18216
rect 6886 18204 6914 18312
rect 10965 18309 10977 18312
rect 11011 18309 11023 18343
rect 10965 18303 11023 18309
rect 17218 18300 17224 18352
rect 17276 18340 17282 18352
rect 17586 18340 17592 18352
rect 17276 18312 17592 18340
rect 17276 18300 17282 18312
rect 17586 18300 17592 18312
rect 17644 18340 17650 18352
rect 18049 18343 18107 18349
rect 18049 18340 18061 18343
rect 17644 18312 18061 18340
rect 17644 18300 17650 18312
rect 18049 18309 18061 18312
rect 18095 18309 18107 18343
rect 32306 18340 32312 18352
rect 32267 18312 32312 18340
rect 18049 18303 18107 18309
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 9122 18272 9128 18284
rect 9083 18244 9128 18272
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18272 17463 18275
rect 17494 18272 17500 18284
rect 17451 18244 17500 18272
rect 17451 18241 17463 18244
rect 17405 18235 17463 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27525 18275 27583 18281
rect 27525 18272 27537 18275
rect 27212 18244 27537 18272
rect 27212 18232 27218 18244
rect 27525 18241 27537 18244
rect 27571 18241 27583 18275
rect 32122 18272 32128 18284
rect 32083 18244 32128 18272
rect 27525 18235 27583 18241
rect 32122 18232 32128 18244
rect 32180 18232 32186 18284
rect 3476 18176 6914 18204
rect 9309 18207 9367 18213
rect 3476 18164 3482 18176
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 33870 18204 33876 18216
rect 33831 18176 33876 18204
rect 9309 18167 9367 18173
rect 6886 18108 8800 18136
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6886 18068 6914 18108
rect 6604 18040 6914 18068
rect 7929 18071 7987 18077
rect 6604 18028 6610 18040
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 8478 18068 8484 18080
rect 7975 18040 8484 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 8662 18068 8668 18080
rect 8623 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8772 18068 8800 18108
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9324 18136 9352 18167
rect 33870 18164 33876 18176
rect 33928 18164 33934 18216
rect 9088 18108 9352 18136
rect 16546 18108 18368 18136
rect 9088 18096 9094 18108
rect 16546 18068 16574 18108
rect 17126 18068 17132 18080
rect 8772 18040 16574 18068
rect 17087 18040 17132 18068
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 18340 18077 18368 18108
rect 18325 18071 18383 18077
rect 18325 18037 18337 18071
rect 18371 18068 18383 18071
rect 27154 18068 27160 18080
rect 18371 18040 27160 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 29546 18068 29552 18080
rect 29507 18040 29552 18068
rect 29546 18028 29552 18040
rect 29604 18028 29610 18080
rect 1104 17978 34868 18000
rect 1104 17926 5174 17978
rect 5226 17926 5238 17978
rect 5290 17926 5302 17978
rect 5354 17926 5366 17978
rect 5418 17926 5430 17978
rect 5482 17926 13622 17978
rect 13674 17926 13686 17978
rect 13738 17926 13750 17978
rect 13802 17926 13814 17978
rect 13866 17926 13878 17978
rect 13930 17926 22070 17978
rect 22122 17926 22134 17978
rect 22186 17926 22198 17978
rect 22250 17926 22262 17978
rect 22314 17926 22326 17978
rect 22378 17926 30518 17978
rect 30570 17926 30582 17978
rect 30634 17926 30646 17978
rect 30698 17926 30710 17978
rect 30762 17926 30774 17978
rect 30826 17926 34868 17978
rect 1104 17904 34868 17926
rect 27249 17867 27307 17873
rect 27249 17833 27261 17867
rect 27295 17864 27307 17867
rect 27338 17864 27344 17876
rect 27295 17836 27344 17864
rect 27295 17833 27307 17836
rect 27249 17827 27307 17833
rect 27338 17824 27344 17836
rect 27396 17824 27402 17876
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 6972 17768 9444 17796
rect 6972 17756 6978 17768
rect 5074 17688 5080 17740
rect 5132 17728 5138 17740
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 5132 17700 5181 17728
rect 5132 17688 5138 17700
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 5169 17691 5227 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 8662 17688 8668 17740
rect 8720 17728 8726 17740
rect 9416 17737 9444 17768
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 8720 17700 8953 17728
rect 8720 17688 8726 17700
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 27798 17688 27804 17740
rect 27856 17728 27862 17740
rect 29546 17728 29552 17740
rect 27856 17700 28856 17728
rect 29507 17700 29552 17728
rect 27856 17688 27862 17700
rect 2038 17660 2044 17672
rect 1999 17632 2044 17660
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 2774 17660 2780 17672
rect 2735 17632 2780 17660
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 17586 17660 17592 17672
rect 17547 17632 17592 17660
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 27154 17660 27160 17672
rect 27115 17632 27160 17660
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 27985 17663 28043 17669
rect 27985 17629 27997 17663
rect 28031 17660 28043 17663
rect 28258 17660 28264 17672
rect 28031 17632 28264 17660
rect 28031 17629 28043 17632
rect 27985 17623 28043 17629
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 28828 17669 28856 17700
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17728 31447 17731
rect 33042 17728 33048 17740
rect 31435 17700 33048 17728
rect 31435 17697 31447 17700
rect 31389 17691 31447 17697
rect 33042 17688 33048 17700
rect 33100 17688 33106 17740
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 5350 17592 5356 17604
rect 5311 17564 5356 17592
rect 5350 17552 5356 17564
rect 5408 17552 5414 17604
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 9125 17595 9183 17601
rect 9125 17592 9137 17595
rect 8536 17564 9137 17592
rect 8536 17552 8542 17564
rect 9125 17561 9137 17564
rect 9171 17561 9183 17595
rect 9125 17555 9183 17561
rect 28905 17595 28963 17601
rect 28905 17561 28917 17595
rect 28951 17592 28963 17595
rect 29733 17595 29791 17601
rect 29733 17592 29745 17595
rect 28951 17564 29745 17592
rect 28951 17561 28963 17564
rect 28905 17555 28963 17561
rect 29733 17561 29745 17564
rect 29779 17561 29791 17595
rect 29733 17555 29791 17561
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1636 17496 1961 17524
rect 1636 17484 1642 17496
rect 1949 17493 1961 17496
rect 1995 17493 2007 17527
rect 1949 17487 2007 17493
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 7834 17524 7840 17536
rect 7432 17496 7840 17524
rect 7432 17484 7438 17496
rect 7834 17484 7840 17496
rect 7892 17524 7898 17536
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 7892 17496 17509 17524
rect 7892 17484 7898 17496
rect 17497 17493 17509 17496
rect 17543 17524 17555 17527
rect 25222 17524 25228 17536
rect 17543 17496 25228 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 27706 17484 27712 17536
rect 27764 17524 27770 17536
rect 27893 17527 27951 17533
rect 27893 17524 27905 17527
rect 27764 17496 27905 17524
rect 27764 17484 27770 17496
rect 27893 17493 27905 17496
rect 27939 17493 27951 17527
rect 27893 17487 27951 17493
rect 1104 17434 34868 17456
rect 1104 17382 9398 17434
rect 9450 17382 9462 17434
rect 9514 17382 9526 17434
rect 9578 17382 9590 17434
rect 9642 17382 9654 17434
rect 9706 17382 17846 17434
rect 17898 17382 17910 17434
rect 17962 17382 17974 17434
rect 18026 17382 18038 17434
rect 18090 17382 18102 17434
rect 18154 17382 26294 17434
rect 26346 17382 26358 17434
rect 26410 17382 26422 17434
rect 26474 17382 26486 17434
rect 26538 17382 26550 17434
rect 26602 17382 34868 17434
rect 1104 17360 34868 17382
rect 2038 17280 2044 17332
rect 2096 17320 2102 17332
rect 5350 17320 5356 17332
rect 2096 17292 3188 17320
rect 5311 17292 5356 17320
rect 2096 17280 2102 17292
rect 3050 17252 3056 17264
rect 2332 17224 3056 17252
rect 2332 17193 2360 17224
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 3160 17252 3188 17292
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 27706 17252 27712 17264
rect 3160 17224 5304 17252
rect 27667 17224 27712 17252
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 2774 17184 2780 17196
rect 2735 17156 2780 17184
rect 2317 17147 2375 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 5276 17193 5304 17224
rect 27706 17212 27712 17224
rect 27764 17212 27770 17264
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2961 17119 3019 17125
rect 2961 17116 2973 17119
rect 2271 17088 2973 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2961 17085 2973 17088
rect 3007 17085 3019 17119
rect 3326 17116 3332 17128
rect 3287 17088 3332 17116
rect 2961 17079 3019 17085
rect 3326 17076 3332 17088
rect 3384 17076 3390 17128
rect 27522 17116 27528 17128
rect 27483 17088 27528 17116
rect 27522 17076 27528 17088
rect 27580 17076 27586 17128
rect 29365 17119 29423 17125
rect 29365 17085 29377 17119
rect 29411 17116 29423 17119
rect 32306 17116 32312 17128
rect 29411 17088 32312 17116
rect 29411 17085 29423 17088
rect 29365 17079 29423 17085
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1489 16983 1547 16989
rect 1489 16980 1501 16983
rect 1452 16952 1501 16980
rect 1452 16940 1458 16952
rect 1489 16949 1501 16952
rect 1535 16949 1547 16983
rect 1489 16943 1547 16949
rect 32306 16940 32312 16992
rect 32364 16980 32370 16992
rect 32861 16983 32919 16989
rect 32861 16980 32873 16983
rect 32364 16952 32873 16980
rect 32364 16940 32370 16952
rect 32861 16949 32873 16952
rect 32907 16949 32919 16983
rect 32861 16943 32919 16949
rect 1104 16890 34868 16912
rect 1104 16838 5174 16890
rect 5226 16838 5238 16890
rect 5290 16838 5302 16890
rect 5354 16838 5366 16890
rect 5418 16838 5430 16890
rect 5482 16838 13622 16890
rect 13674 16838 13686 16890
rect 13738 16838 13750 16890
rect 13802 16838 13814 16890
rect 13866 16838 13878 16890
rect 13930 16838 22070 16890
rect 22122 16838 22134 16890
rect 22186 16838 22198 16890
rect 22250 16838 22262 16890
rect 22314 16838 22326 16890
rect 22378 16838 30518 16890
rect 30570 16838 30582 16890
rect 30634 16838 30646 16890
rect 30698 16838 30710 16890
rect 30762 16838 30774 16890
rect 30826 16838 34868 16890
rect 1104 16816 34868 16838
rect 27522 16736 27528 16788
rect 27580 16776 27586 16788
rect 27617 16779 27675 16785
rect 27617 16776 27629 16779
rect 27580 16748 27629 16776
rect 27580 16736 27586 16748
rect 27617 16745 27629 16748
rect 27663 16745 27675 16779
rect 27617 16739 27675 16745
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 32306 16640 32312 16652
rect 32267 16612 32312 16640
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 3234 16572 3240 16584
rect 3195 16544 3240 16572
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 32493 16507 32551 16513
rect 32493 16473 32505 16507
rect 32539 16504 32551 16507
rect 32766 16504 32772 16516
rect 32539 16476 32772 16504
rect 32539 16473 32551 16476
rect 32493 16467 32551 16473
rect 32766 16464 32772 16476
rect 32824 16464 32830 16516
rect 34146 16504 34152 16516
rect 34107 16476 34152 16504
rect 34146 16464 34152 16476
rect 34204 16464 34210 16516
rect 1104 16346 34868 16368
rect 1104 16294 9398 16346
rect 9450 16294 9462 16346
rect 9514 16294 9526 16346
rect 9578 16294 9590 16346
rect 9642 16294 9654 16346
rect 9706 16294 17846 16346
rect 17898 16294 17910 16346
rect 17962 16294 17974 16346
rect 18026 16294 18038 16346
rect 18090 16294 18102 16346
rect 18154 16294 26294 16346
rect 26346 16294 26358 16346
rect 26410 16294 26422 16346
rect 26474 16294 26486 16346
rect 26538 16294 26550 16346
rect 26602 16294 34868 16346
rect 1104 16272 34868 16294
rect 32766 16232 32772 16244
rect 32727 16204 32772 16232
rect 32766 16192 32772 16204
rect 32824 16192 32830 16244
rect 17402 16164 17408 16176
rect 17363 16136 17408 16164
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 18230 16124 18236 16176
rect 18288 16164 18294 16176
rect 33134 16164 33140 16176
rect 18288 16136 33140 16164
rect 18288 16124 18294 16136
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 18248 16096 18276 16124
rect 32876 16105 32904 16136
rect 33134 16124 33140 16136
rect 33192 16124 33198 16176
rect 9171 16068 18276 16096
rect 32861 16099 32919 16105
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 32861 16065 32873 16099
rect 32907 16065 32919 16099
rect 32861 16059 32919 16065
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 16028 21327 16031
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21315 16000 21833 16028
rect 21315 15997 21327 16000
rect 21269 15991 21327 15997
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 23661 16031 23719 16037
rect 23661 15997 23673 16031
rect 23707 16028 23719 16031
rect 32398 16028 32404 16040
rect 23707 16000 32404 16028
rect 23707 15997 23719 16000
rect 23661 15991 23719 15997
rect 20806 15920 20812 15972
rect 20864 15960 20870 15972
rect 22020 15960 22048 15991
rect 32398 15988 32404 16000
rect 32456 15988 32462 16040
rect 20864 15932 22048 15960
rect 20864 15920 20870 15932
rect 4246 15892 4252 15904
rect 4207 15864 4252 15892
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 8938 15892 8944 15904
rect 8527 15864 8944 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9033 15895 9091 15901
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 9122 15892 9128 15904
rect 9079 15864 9128 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17129 15895 17187 15901
rect 17129 15892 17141 15895
rect 17000 15864 17141 15892
rect 17000 15852 17006 15864
rect 17129 15861 17141 15864
rect 17175 15861 17187 15895
rect 17129 15855 17187 15861
rect 1104 15802 34868 15824
rect 1104 15750 5174 15802
rect 5226 15750 5238 15802
rect 5290 15750 5302 15802
rect 5354 15750 5366 15802
rect 5418 15750 5430 15802
rect 5482 15750 13622 15802
rect 13674 15750 13686 15802
rect 13738 15750 13750 15802
rect 13802 15750 13814 15802
rect 13866 15750 13878 15802
rect 13930 15750 22070 15802
rect 22122 15750 22134 15802
rect 22186 15750 22198 15802
rect 22250 15750 22262 15802
rect 22314 15750 22326 15802
rect 22378 15750 30518 15802
rect 30570 15750 30582 15802
rect 30634 15750 30646 15802
rect 30698 15750 30710 15802
rect 30762 15750 30774 15802
rect 30826 15750 34868 15802
rect 1104 15728 34868 15750
rect 20806 15688 20812 15700
rect 20767 15660 20812 15688
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 4062 15580 4068 15632
rect 4120 15620 4126 15632
rect 4120 15592 4752 15620
rect 4120 15580 4126 15592
rect 4246 15552 4252 15564
rect 4207 15524 4252 15552
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4724 15561 4752 15592
rect 4709 15555 4767 15561
rect 4709 15521 4721 15555
rect 4755 15521 4767 15555
rect 8938 15552 8944 15564
rect 8899 15524 8944 15552
rect 4709 15515 4767 15521
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9122 15552 9128 15564
rect 9083 15524 9128 15552
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 9858 15552 9864 15564
rect 9819 15524 9864 15552
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 17402 15444 17408 15496
rect 17460 15484 17466 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17460 15456 17693 15484
rect 17460 15444 17466 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 20717 15487 20775 15493
rect 20717 15484 20729 15487
rect 19024 15456 20729 15484
rect 19024 15444 19030 15456
rect 20717 15453 20729 15456
rect 20763 15484 20775 15487
rect 20990 15484 20996 15496
rect 20763 15456 20996 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 4430 15416 4436 15428
rect 4391 15388 4436 15416
rect 4430 15376 4436 15388
rect 4488 15376 4494 15428
rect 17494 15348 17500 15360
rect 17407 15320 17500 15348
rect 17494 15308 17500 15320
rect 17552 15348 17558 15360
rect 18966 15348 18972 15360
rect 17552 15320 18972 15348
rect 17552 15308 17558 15320
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 1104 15258 34868 15280
rect 1104 15206 9398 15258
rect 9450 15206 9462 15258
rect 9514 15206 9526 15258
rect 9578 15206 9590 15258
rect 9642 15206 9654 15258
rect 9706 15206 17846 15258
rect 17898 15206 17910 15258
rect 17962 15206 17974 15258
rect 18026 15206 18038 15258
rect 18090 15206 18102 15258
rect 18154 15206 26294 15258
rect 26346 15206 26358 15258
rect 26410 15206 26422 15258
rect 26474 15206 26486 15258
rect 26538 15206 26550 15258
rect 26602 15206 34868 15258
rect 1104 15184 34868 15206
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 4488 15116 4813 15144
rect 4488 15104 4494 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 4801 15107 4859 15113
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 17494 15144 17500 15156
rect 10284 15116 17500 15144
rect 10284 15104 10290 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 1946 15008 1952 15020
rect 1907 14980 1952 15008
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5626 15008 5632 15020
rect 4939 14980 5632 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 15008 18935 15011
rect 18966 15008 18972 15020
rect 18923 14980 18972 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 25225 15011 25283 15017
rect 25225 14977 25237 15011
rect 25271 15008 25283 15011
rect 27154 15008 27160 15020
rect 25271 14980 27160 15008
rect 25271 14977 25283 14980
rect 25225 14971 25283 14977
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 19150 14940 19156 14952
rect 19063 14912 19156 14940
rect 19150 14900 19156 14912
rect 19208 14940 19214 14952
rect 31018 14940 31024 14952
rect 19208 14912 31024 14940
rect 19208 14900 19214 14912
rect 31018 14900 31024 14912
rect 31076 14940 31082 14952
rect 31938 14940 31944 14952
rect 31076 14912 31944 14940
rect 31076 14900 31082 14912
rect 31938 14900 31944 14912
rect 31996 14900 32002 14952
rect 1578 14764 1584 14816
rect 1636 14804 1642 14816
rect 1857 14807 1915 14813
rect 1857 14804 1869 14807
rect 1636 14776 1869 14804
rect 1636 14764 1642 14776
rect 1857 14773 1869 14776
rect 1903 14773 1915 14807
rect 1857 14767 1915 14773
rect 25317 14807 25375 14813
rect 25317 14773 25329 14807
rect 25363 14804 25375 14807
rect 25498 14804 25504 14816
rect 25363 14776 25504 14804
rect 25363 14773 25375 14776
rect 25317 14767 25375 14773
rect 25498 14764 25504 14776
rect 25556 14764 25562 14816
rect 1104 14714 34868 14736
rect 1104 14662 5174 14714
rect 5226 14662 5238 14714
rect 5290 14662 5302 14714
rect 5354 14662 5366 14714
rect 5418 14662 5430 14714
rect 5482 14662 13622 14714
rect 13674 14662 13686 14714
rect 13738 14662 13750 14714
rect 13802 14662 13814 14714
rect 13866 14662 13878 14714
rect 13930 14662 22070 14714
rect 22122 14662 22134 14714
rect 22186 14662 22198 14714
rect 22250 14662 22262 14714
rect 22314 14662 22326 14714
rect 22378 14662 30518 14714
rect 30570 14662 30582 14714
rect 30634 14662 30646 14714
rect 30698 14662 30710 14714
rect 30762 14662 30774 14714
rect 30826 14662 34868 14714
rect 1104 14640 34868 14662
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 1854 14464 1860 14476
rect 1815 14436 1860 14464
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 25498 14464 25504 14476
rect 25459 14436 25504 14464
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 25314 14396 25320 14408
rect 25275 14368 25320 14396
rect 25314 14356 25320 14368
rect 25372 14356 25378 14408
rect 27157 14331 27215 14337
rect 27157 14297 27169 14331
rect 27203 14328 27215 14331
rect 31754 14328 31760 14340
rect 27203 14300 31760 14328
rect 27203 14297 27215 14300
rect 27157 14291 27215 14297
rect 31754 14288 31760 14300
rect 31812 14288 31818 14340
rect 1104 14170 34868 14192
rect 1104 14118 9398 14170
rect 9450 14118 9462 14170
rect 9514 14118 9526 14170
rect 9578 14118 9590 14170
rect 9642 14118 9654 14170
rect 9706 14118 17846 14170
rect 17898 14118 17910 14170
rect 17962 14118 17974 14170
rect 18026 14118 18038 14170
rect 18090 14118 18102 14170
rect 18154 14118 26294 14170
rect 26346 14118 26358 14170
rect 26410 14118 26422 14170
rect 26474 14118 26486 14170
rect 26538 14118 26550 14170
rect 26602 14118 34868 14170
rect 1104 14096 34868 14118
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1489 13923 1547 13929
rect 1489 13920 1501 13923
rect 1452 13892 1501 13920
rect 1452 13880 1458 13892
rect 1489 13889 1501 13892
rect 1535 13889 1547 13923
rect 6546 13920 6552 13932
rect 6507 13892 6552 13920
rect 1489 13883 1547 13889
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 17678 13920 17684 13932
rect 17639 13892 17684 13920
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 25314 13920 25320 13932
rect 25275 13892 25320 13920
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 6178 13852 6184 13864
rect 5491 13824 6184 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6457 13855 6515 13861
rect 6457 13821 6469 13855
rect 6503 13852 6515 13855
rect 6914 13852 6920 13864
rect 6503 13824 6920 13852
rect 6503 13821 6515 13824
rect 6457 13815 6515 13821
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 16850 13716 16856 13728
rect 16811 13688 16856 13716
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 17589 13719 17647 13725
rect 17589 13716 17601 13719
rect 17092 13688 17601 13716
rect 17092 13676 17098 13688
rect 17589 13685 17601 13688
rect 17635 13685 17647 13719
rect 25958 13716 25964 13728
rect 25919 13688 25964 13716
rect 17589 13679 17647 13685
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 32306 13676 32312 13728
rect 32364 13716 32370 13728
rect 32769 13719 32827 13725
rect 32769 13716 32781 13719
rect 32364 13688 32781 13716
rect 32364 13676 32370 13688
rect 32769 13685 32781 13688
rect 32815 13685 32827 13719
rect 33962 13716 33968 13728
rect 33923 13688 33968 13716
rect 32769 13679 32827 13685
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 1104 13626 34868 13648
rect 1104 13574 5174 13626
rect 5226 13574 5238 13626
rect 5290 13574 5302 13626
rect 5354 13574 5366 13626
rect 5418 13574 5430 13626
rect 5482 13574 13622 13626
rect 13674 13574 13686 13626
rect 13738 13574 13750 13626
rect 13802 13574 13814 13626
rect 13866 13574 13878 13626
rect 13930 13574 22070 13626
rect 22122 13574 22134 13626
rect 22186 13574 22198 13626
rect 22250 13574 22262 13626
rect 22314 13574 22326 13626
rect 22378 13574 30518 13626
rect 30570 13574 30582 13626
rect 30634 13574 30646 13626
rect 30698 13574 30710 13626
rect 30762 13574 30774 13626
rect 30826 13574 34868 13626
rect 1104 13552 34868 13574
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 6236 13416 6914 13444
rect 6236 13404 6242 13416
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 2832 13348 5273 13376
rect 2832 13336 2838 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 6886 13376 6914 13416
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 16816 13416 17356 13444
rect 16816 13404 16822 13416
rect 7101 13379 7159 13385
rect 7101 13376 7113 13379
rect 6886 13348 7113 13376
rect 5261 13339 5319 13345
rect 7101 13345 7113 13348
rect 7147 13345 7159 13379
rect 16850 13376 16856 13388
rect 16811 13348 16856 13376
rect 7101 13339 7159 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 17034 13376 17040 13388
rect 16995 13348 17040 13376
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 17328 13385 17356 13416
rect 17313 13379 17371 13385
rect 17313 13345 17325 13379
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 25409 13379 25467 13385
rect 25409 13345 25421 13379
rect 25455 13376 25467 13379
rect 25958 13376 25964 13388
rect 25455 13348 25964 13376
rect 25455 13345 25467 13348
rect 25409 13339 25467 13345
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 27249 13379 27307 13385
rect 27249 13345 27261 13379
rect 27295 13376 27307 13379
rect 32766 13376 32772 13388
rect 27295 13348 32772 13376
rect 27295 13345 27307 13348
rect 27249 13339 27307 13345
rect 32766 13336 32772 13348
rect 32824 13336 32830 13388
rect 33042 13376 33048 13388
rect 33003 13348 33048 13376
rect 33042 13336 33048 13348
rect 33100 13336 33106 13388
rect 33962 13336 33968 13388
rect 34020 13376 34026 13388
rect 34149 13379 34207 13385
rect 34149 13376 34161 13379
rect 34020 13348 34161 13376
rect 34020 13336 34026 13348
rect 34149 13345 34161 13348
rect 34195 13345 34207 13379
rect 34149 13339 34207 13345
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13308 7803 13311
rect 8202 13308 8208 13320
rect 7791 13280 8208 13308
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10226 13308 10232 13320
rect 10008 13280 10232 13308
rect 10008 13268 10014 13280
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 25590 13240 25596 13252
rect 6972 13212 7017 13240
rect 25551 13212 25596 13240
rect 6972 13200 6978 13212
rect 25590 13200 25596 13212
rect 25648 13200 25654 13252
rect 33962 13240 33968 13252
rect 33923 13212 33968 13240
rect 33962 13200 33968 13212
rect 34020 13200 34026 13252
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 1104 13082 34868 13104
rect 1104 13030 9398 13082
rect 9450 13030 9462 13082
rect 9514 13030 9526 13082
rect 9578 13030 9590 13082
rect 9642 13030 9654 13082
rect 9706 13030 17846 13082
rect 17898 13030 17910 13082
rect 17962 13030 17974 13082
rect 18026 13030 18038 13082
rect 18090 13030 18102 13082
rect 18154 13030 26294 13082
rect 26346 13030 26358 13082
rect 26410 13030 26422 13082
rect 26474 13030 26486 13082
rect 26538 13030 26550 13082
rect 26602 13030 34868 13082
rect 1104 13008 34868 13030
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 14366 12968 14372 12980
rect 5684 12940 14372 12968
rect 5684 12928 5690 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 25409 12971 25467 12977
rect 25409 12937 25421 12971
rect 25455 12968 25467 12971
rect 25590 12968 25596 12980
rect 25455 12940 25596 12968
rect 25455 12937 25467 12940
rect 25409 12931 25467 12937
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 5721 12903 5779 12909
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 8021 12903 8079 12909
rect 8021 12900 8033 12903
rect 5767 12872 8033 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 8021 12869 8033 12872
rect 8067 12869 8079 12903
rect 34146 12900 34152 12912
rect 34107 12872 34152 12900
rect 8021 12863 8079 12869
rect 34146 12860 34152 12872
rect 34204 12860 34210 12912
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 25314 12832 25320 12844
rect 8260 12804 8305 12832
rect 25275 12804 25320 12832
rect 8260 12792 8266 12804
rect 25314 12792 25320 12804
rect 25372 12792 25378 12844
rect 32306 12832 32312 12844
rect 32267 12804 32312 12832
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 6365 12767 6423 12773
rect 6365 12764 6377 12767
rect 4212 12736 6377 12764
rect 4212 12724 4218 12736
rect 6365 12733 6377 12736
rect 6411 12733 6423 12767
rect 32490 12764 32496 12776
rect 32451 12736 32496 12764
rect 6365 12727 6423 12733
rect 32490 12724 32496 12736
rect 32548 12724 32554 12776
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 16298 12628 16304 12640
rect 14424 12600 16304 12628
rect 14424 12588 14430 12600
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 1104 12538 34868 12560
rect 1104 12486 5174 12538
rect 5226 12486 5238 12538
rect 5290 12486 5302 12538
rect 5354 12486 5366 12538
rect 5418 12486 5430 12538
rect 5482 12486 13622 12538
rect 13674 12486 13686 12538
rect 13738 12486 13750 12538
rect 13802 12486 13814 12538
rect 13866 12486 13878 12538
rect 13930 12486 22070 12538
rect 22122 12486 22134 12538
rect 22186 12486 22198 12538
rect 22250 12486 22262 12538
rect 22314 12486 22326 12538
rect 22378 12486 30518 12538
rect 30570 12486 30582 12538
rect 30634 12486 30646 12538
rect 30698 12486 30710 12538
rect 30762 12486 30774 12538
rect 30826 12486 34868 12538
rect 1104 12464 34868 12486
rect 32490 12384 32496 12436
rect 32548 12424 32554 12436
rect 32585 12427 32643 12433
rect 32585 12424 32597 12427
rect 32548 12396 32597 12424
rect 32548 12384 32554 12396
rect 32585 12393 32597 12396
rect 32631 12393 32643 12427
rect 32585 12387 32643 12393
rect 33873 12427 33931 12433
rect 33873 12393 33885 12427
rect 33919 12424 33931 12427
rect 33962 12424 33968 12436
rect 33919 12396 33968 12424
rect 33919 12393 33931 12396
rect 33873 12387 33931 12393
rect 33962 12384 33968 12396
rect 34020 12384 34026 12436
rect 32490 12220 32496 12232
rect 32451 12192 32496 12220
rect 32490 12180 32496 12192
rect 32548 12180 32554 12232
rect 33778 12220 33784 12232
rect 33739 12192 33784 12220
rect 33778 12180 33784 12192
rect 33836 12180 33842 12232
rect 1104 11994 34868 12016
rect 1104 11942 9398 11994
rect 9450 11942 9462 11994
rect 9514 11942 9526 11994
rect 9578 11942 9590 11994
rect 9642 11942 9654 11994
rect 9706 11942 17846 11994
rect 17898 11942 17910 11994
rect 17962 11942 17974 11994
rect 18026 11942 18038 11994
rect 18090 11942 18102 11994
rect 18154 11942 26294 11994
rect 26346 11942 26358 11994
rect 26410 11942 26422 11994
rect 26474 11942 26486 11994
rect 26538 11942 26550 11994
rect 26602 11942 34868 11994
rect 1104 11920 34868 11942
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17770 11744 17776 11756
rect 17635 11716 17776 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20806 11744 20812 11756
rect 20763 11716 20812 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 14274 11540 14280 11552
rect 14235 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16908 11512 16957 11540
rect 16908 11500 16914 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17497 11543 17555 11549
rect 17497 11540 17509 11543
rect 17092 11512 17509 11540
rect 17092 11500 17098 11512
rect 17497 11509 17509 11512
rect 17543 11509 17555 11543
rect 17497 11503 17555 11509
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 20898 11540 20904 11552
rect 20855 11512 20904 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 34868 11472
rect 1104 11398 5174 11450
rect 5226 11398 5238 11450
rect 5290 11398 5302 11450
rect 5354 11398 5366 11450
rect 5418 11398 5430 11450
rect 5482 11398 13622 11450
rect 13674 11398 13686 11450
rect 13738 11398 13750 11450
rect 13802 11398 13814 11450
rect 13866 11398 13878 11450
rect 13930 11398 22070 11450
rect 22122 11398 22134 11450
rect 22186 11398 22198 11450
rect 22250 11398 22262 11450
rect 22314 11398 22326 11450
rect 22378 11398 30518 11450
rect 30570 11398 30582 11450
rect 30634 11398 30646 11450
rect 30698 11398 30710 11450
rect 30762 11398 30774 11450
rect 30826 11398 34868 11450
rect 1104 11376 34868 11398
rect 6886 11240 17356 11268
rect 658 11160 664 11212
rect 716 11200 722 11212
rect 6886 11200 6914 11240
rect 14274 11200 14280 11212
rect 716 11172 6914 11200
rect 14235 11172 14280 11200
rect 716 11160 722 11172
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14826 11200 14832 11212
rect 14787 11172 14832 11200
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 16850 11200 16856 11212
rect 16811 11172 16856 11200
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 17034 11200 17040 11212
rect 16995 11172 17040 11200
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17328 11209 17356 11240
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11169 17371 11203
rect 20898 11200 20904 11212
rect 20859 11172 20904 11200
rect 17313 11163 17371 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 21726 11200 21732 11212
rect 21687 11172 21732 11200
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7340 11104 7385 11132
rect 7340 11092 7346 11104
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 9180 11104 9229 11132
rect 9180 11092 9186 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 20714 11132 20720 11144
rect 20675 11104 20720 11132
rect 9217 11095 9275 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 5445 11067 5503 11073
rect 5445 11064 5457 11067
rect 3384 11036 5457 11064
rect 3384 11024 3390 11036
rect 5445 11033 5457 11036
rect 5491 11033 5503 11067
rect 7098 11064 7104 11076
rect 7059 11036 7104 11064
rect 5445 11027 5503 11033
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 14458 11064 14464 11076
rect 14419 11036 14464 11064
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 2866 10996 2872 11008
rect 2827 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 1104 10906 34868 10928
rect 1104 10854 9398 10906
rect 9450 10854 9462 10906
rect 9514 10854 9526 10906
rect 9578 10854 9590 10906
rect 9642 10854 9654 10906
rect 9706 10854 17846 10906
rect 17898 10854 17910 10906
rect 17962 10854 17974 10906
rect 18026 10854 18038 10906
rect 18090 10854 18102 10906
rect 18154 10854 26294 10906
rect 26346 10854 26358 10906
rect 26410 10854 26422 10906
rect 26474 10854 26486 10906
rect 26538 10854 26550 10906
rect 26602 10854 34868 10906
rect 1104 10832 34868 10854
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 7098 10792 7104 10804
rect 6503 10764 7104 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 14458 10792 14464 10804
rect 14419 10764 14464 10792
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 2866 10724 2872 10736
rect 2639 10696 2872 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 17678 10724 17684 10736
rect 6886 10696 17684 10724
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 2372 10628 2421 10656
rect 2372 10616 2378 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6886 10656 6914 10696
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 27249 10727 27307 10733
rect 27249 10693 27261 10727
rect 27295 10724 27307 10727
rect 27985 10727 28043 10733
rect 27985 10724 27997 10727
rect 27295 10696 27997 10724
rect 27295 10693 27307 10696
rect 27249 10687 27307 10693
rect 27985 10693 27997 10696
rect 28031 10693 28043 10727
rect 27985 10687 28043 10693
rect 9122 10656 9128 10668
rect 6595 10628 6914 10656
rect 9083 10628 9128 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 14366 10656 14372 10668
rect 14327 10628 14372 10656
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27120 10628 27169 10656
rect 27120 10616 27126 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2832 10560 2881 10588
rect 2832 10548 2838 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 7282 10588 7288 10600
rect 5767 10560 7288 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9766 10588 9772 10600
rect 9355 10560 9772 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 27798 10588 27804 10600
rect 27759 10560 27804 10588
rect 9861 10551 9919 10557
rect 8938 10480 8944 10532
rect 8996 10520 9002 10532
rect 9876 10520 9904 10551
rect 27798 10548 27804 10560
rect 27856 10548 27862 10600
rect 29641 10591 29699 10597
rect 29641 10557 29653 10591
rect 29687 10588 29699 10591
rect 31662 10588 31668 10600
rect 29687 10560 31668 10588
rect 29687 10557 29699 10560
rect 29641 10551 29699 10557
rect 31662 10548 31668 10560
rect 31720 10548 31726 10600
rect 8996 10492 9904 10520
rect 8996 10480 9002 10492
rect 1104 10362 34868 10384
rect 1104 10310 5174 10362
rect 5226 10310 5238 10362
rect 5290 10310 5302 10362
rect 5354 10310 5366 10362
rect 5418 10310 5430 10362
rect 5482 10310 13622 10362
rect 13674 10310 13686 10362
rect 13738 10310 13750 10362
rect 13802 10310 13814 10362
rect 13866 10310 13878 10362
rect 13930 10310 22070 10362
rect 22122 10310 22134 10362
rect 22186 10310 22198 10362
rect 22250 10310 22262 10362
rect 22314 10310 22326 10362
rect 22378 10310 30518 10362
rect 30570 10310 30582 10362
rect 30634 10310 30646 10362
rect 30698 10310 30710 10362
rect 30762 10310 30774 10362
rect 30826 10310 34868 10362
rect 1104 10288 34868 10310
rect 9766 10248 9772 10260
rect 9727 10220 9772 10248
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 27798 10208 27804 10260
rect 27856 10248 27862 10260
rect 27893 10251 27951 10257
rect 27893 10248 27905 10251
rect 27856 10220 27905 10248
rect 27856 10208 27862 10220
rect 27893 10217 27905 10220
rect 27939 10217 27951 10251
rect 27893 10211 27951 10217
rect 1946 10112 1952 10124
rect 1780 10084 1952 10112
rect 1780 10053 1808 10084
rect 1946 10072 1952 10084
rect 2004 10112 2010 10124
rect 10410 10112 10416 10124
rect 2004 10084 10416 10112
rect 2004 10072 2010 10084
rect 10410 10072 10416 10084
rect 10468 10112 10474 10124
rect 10468 10084 11376 10112
rect 10468 10072 10474 10084
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 1765 10007 1823 10013
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 11348 10053 11376 10084
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 3016 10016 3065 10044
rect 3016 10004 3022 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 9876 9976 9904 10007
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11940 10016 11989 10044
rect 11940 10004 11946 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 19521 10047 19579 10053
rect 19521 10044 19533 10047
rect 16540 10016 19533 10044
rect 16540 10004 16546 10016
rect 19521 10013 19533 10016
rect 19567 10044 19579 10047
rect 28258 10044 28264 10056
rect 19567 10016 28264 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 12158 9976 12164 9988
rect 9876 9948 12164 9976
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 1673 9911 1731 9917
rect 1673 9908 1685 9911
rect 1636 9880 1685 9908
rect 1636 9868 1642 9880
rect 1673 9877 1685 9880
rect 1719 9877 1731 9911
rect 2958 9908 2964 9920
rect 2919 9880 2964 9908
rect 1673 9871 1731 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 11425 9911 11483 9917
rect 11425 9877 11437 9911
rect 11471 9908 11483 9911
rect 12066 9908 12072 9920
rect 11471 9880 12072 9908
rect 11471 9877 11483 9880
rect 11425 9871 11483 9877
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 16666 9908 16672 9920
rect 16540 9880 16672 9908
rect 16540 9868 16546 9880
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 19610 9908 19616 9920
rect 19571 9880 19616 9908
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 1104 9818 34868 9840
rect 1104 9766 9398 9818
rect 9450 9766 9462 9818
rect 9514 9766 9526 9818
rect 9578 9766 9590 9818
rect 9642 9766 9654 9818
rect 9706 9766 17846 9818
rect 17898 9766 17910 9818
rect 17962 9766 17974 9818
rect 18026 9766 18038 9818
rect 18090 9766 18102 9818
rect 18154 9766 26294 9818
rect 26346 9766 26358 9818
rect 26410 9766 26422 9818
rect 26474 9766 26486 9818
rect 26538 9766 26550 9818
rect 26602 9766 34868 9818
rect 1104 9744 34868 9766
rect 2685 9639 2743 9645
rect 2685 9605 2697 9639
rect 2731 9636 2743 9639
rect 2958 9636 2964 9648
rect 2731 9608 2964 9636
rect 2731 9605 2743 9608
rect 2685 9599 2743 9605
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 12066 9636 12072 9648
rect 12027 9608 12072 9636
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 12158 9596 12164 9648
rect 12216 9636 12222 9648
rect 16482 9636 16488 9648
rect 12216 9608 16488 9636
rect 12216 9596 12222 9608
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 19610 9636 19616 9648
rect 19571 9608 19616 9636
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2464 9540 2513 9568
rect 2464 9528 2470 9540
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 11882 9568 11888 9580
rect 11843 9540 11888 9568
rect 2501 9531 2559 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 2832 9472 2973 9500
rect 2832 9460 2838 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 13446 9500 13452 9512
rect 13407 9472 13452 9500
rect 2961 9463 3019 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 19426 9500 19432 9512
rect 19387 9472 19432 9500
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19978 9500 19984 9512
rect 19939 9472 19984 9500
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1489 9367 1547 9373
rect 1489 9364 1501 9367
rect 1452 9336 1501 9364
rect 1452 9324 1458 9336
rect 1489 9333 1501 9336
rect 1535 9333 1547 9367
rect 1489 9327 1547 9333
rect 1104 9274 34868 9296
rect 1104 9222 5174 9274
rect 5226 9222 5238 9274
rect 5290 9222 5302 9274
rect 5354 9222 5366 9274
rect 5418 9222 5430 9274
rect 5482 9222 13622 9274
rect 13674 9222 13686 9274
rect 13738 9222 13750 9274
rect 13802 9222 13814 9274
rect 13866 9222 13878 9274
rect 13930 9222 22070 9274
rect 22122 9222 22134 9274
rect 22186 9222 22198 9274
rect 22250 9222 22262 9274
rect 22314 9222 22326 9274
rect 22378 9222 30518 9274
rect 30570 9222 30582 9274
rect 30634 9222 30646 9274
rect 30698 9222 30710 9274
rect 30762 9222 30774 9274
rect 30826 9222 34868 9274
rect 1104 9200 34868 9222
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19521 9163 19579 9169
rect 19521 9160 19533 9163
rect 19484 9132 19533 9160
rect 19484 9120 19490 9132
rect 19521 9129 19533 9132
rect 19567 9129 19579 9163
rect 19521 9123 19579 9129
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 8984 1458 9036
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 1854 9024 1860 9036
rect 1815 8996 1860 9024
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 20864 8996 24624 9024
rect 20864 8984 20870 8996
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 23934 8956 23940 8968
rect 23891 8928 23940 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 24596 8965 24624 8996
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 30926 8956 30932 8968
rect 30887 8928 30932 8956
rect 24581 8919 24639 8925
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 30834 8848 30840 8900
rect 30892 8888 30898 8900
rect 31113 8891 31171 8897
rect 31113 8888 31125 8891
rect 30892 8860 31125 8888
rect 30892 8848 30898 8860
rect 31113 8857 31125 8860
rect 31159 8857 31171 8891
rect 32766 8888 32772 8900
rect 32727 8860 32772 8888
rect 31113 8851 31171 8857
rect 32766 8848 32772 8860
rect 32824 8848 32830 8900
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 24176 8792 24501 8820
rect 24176 8780 24182 8792
rect 24489 8789 24501 8792
rect 24535 8789 24547 8823
rect 24489 8783 24547 8789
rect 1104 8730 34868 8752
rect 1104 8678 9398 8730
rect 9450 8678 9462 8730
rect 9514 8678 9526 8730
rect 9578 8678 9590 8730
rect 9642 8678 9654 8730
rect 9706 8678 17846 8730
rect 17898 8678 17910 8730
rect 17962 8678 17974 8730
rect 18026 8678 18038 8730
rect 18090 8678 18102 8730
rect 18154 8678 26294 8730
rect 26346 8678 26358 8730
rect 26410 8678 26422 8730
rect 26474 8678 26486 8730
rect 26538 8678 26550 8730
rect 26602 8678 34868 8730
rect 1104 8656 34868 8678
rect 30834 8616 30840 8628
rect 30795 8588 30840 8616
rect 30834 8576 30840 8588
rect 30892 8576 30898 8628
rect 24118 8548 24124 8560
rect 24079 8520 24124 8548
rect 24118 8508 24124 8520
rect 24176 8508 24182 8560
rect 31018 8548 31024 8560
rect 30760 8520 31024 8548
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 12158 8480 12164 8492
rect 11747 8452 12164 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 23934 8480 23940 8492
rect 23895 8452 23940 8480
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 28258 8440 28264 8492
rect 28316 8480 28322 8492
rect 30760 8489 30788 8520
rect 31018 8508 31024 8520
rect 31076 8508 31082 8560
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28316 8452 29101 8480
rect 28316 8440 28322 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 30745 8483 30803 8489
rect 30745 8449 30757 8483
rect 30791 8449 30803 8483
rect 30745 8443 30803 8449
rect 30926 8440 30932 8492
rect 30984 8480 30990 8492
rect 31389 8483 31447 8489
rect 31389 8480 31401 8483
rect 30984 8452 31401 8480
rect 30984 8440 30990 8452
rect 31389 8449 31401 8452
rect 31435 8449 31447 8483
rect 31389 8443 31447 8449
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8412 11667 8415
rect 12894 8412 12900 8424
rect 11655 8384 12900 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 24486 8412 24492 8424
rect 24447 8384 24492 8412
rect 24486 8372 24492 8384
rect 24544 8372 24550 8424
rect 12345 8347 12403 8353
rect 12345 8313 12357 8347
rect 12391 8344 12403 8347
rect 13078 8344 13084 8356
rect 12391 8316 13084 8344
rect 12391 8313 12403 8316
rect 12345 8307 12403 8313
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 9858 8276 9864 8288
rect 3200 8248 9864 8276
rect 3200 8236 3206 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 29178 8276 29184 8288
rect 29139 8248 29184 8276
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 29730 8276 29736 8288
rect 29691 8248 29736 8276
rect 29730 8236 29736 8248
rect 29788 8236 29794 8288
rect 1104 8186 34868 8208
rect 1104 8134 5174 8186
rect 5226 8134 5238 8186
rect 5290 8134 5302 8186
rect 5354 8134 5366 8186
rect 5418 8134 5430 8186
rect 5482 8134 13622 8186
rect 13674 8134 13686 8186
rect 13738 8134 13750 8186
rect 13802 8134 13814 8186
rect 13866 8134 13878 8186
rect 13930 8134 22070 8186
rect 22122 8134 22134 8186
rect 22186 8134 22198 8186
rect 22250 8134 22262 8186
rect 22314 8134 22326 8186
rect 22378 8134 30518 8186
rect 30570 8134 30582 8186
rect 30634 8134 30646 8186
rect 30698 8134 30710 8186
rect 30762 8134 30774 8186
rect 30826 8134 34868 8186
rect 1104 8112 34868 8134
rect 12894 7936 12900 7948
rect 12855 7908 12900 7936
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 13078 7936 13084 7948
rect 13039 7908 13084 7936
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 29549 7939 29607 7945
rect 29549 7905 29561 7939
rect 29595 7936 29607 7939
rect 29730 7936 29736 7948
rect 29595 7908 29736 7936
rect 29595 7905 29607 7908
rect 29549 7899 29607 7905
rect 29730 7896 29736 7908
rect 29788 7896 29794 7948
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 11241 7803 11299 7809
rect 11241 7800 11253 7803
rect 10100 7772 11253 7800
rect 10100 7760 10106 7772
rect 11241 7769 11253 7772
rect 11287 7769 11299 7803
rect 11241 7763 11299 7769
rect 29178 7760 29184 7812
rect 29236 7800 29242 7812
rect 29733 7803 29791 7809
rect 29733 7800 29745 7803
rect 29236 7772 29745 7800
rect 29236 7760 29242 7772
rect 29733 7769 29745 7772
rect 29779 7769 29791 7803
rect 29733 7763 29791 7769
rect 31389 7803 31447 7809
rect 31389 7769 31401 7803
rect 31435 7800 31447 7803
rect 33042 7800 33048 7812
rect 31435 7772 33048 7800
rect 31435 7769 31447 7772
rect 31389 7763 31447 7769
rect 33042 7760 33048 7772
rect 33100 7760 33106 7812
rect 1104 7642 34868 7664
rect 1104 7590 9398 7642
rect 9450 7590 9462 7642
rect 9514 7590 9526 7642
rect 9578 7590 9590 7642
rect 9642 7590 9654 7642
rect 9706 7590 17846 7642
rect 17898 7590 17910 7642
rect 17962 7590 17974 7642
rect 18026 7590 18038 7642
rect 18090 7590 18102 7642
rect 18154 7590 26294 7642
rect 26346 7590 26358 7642
rect 26410 7590 26422 7642
rect 26474 7590 26486 7642
rect 26538 7590 26550 7642
rect 26602 7590 34868 7642
rect 1104 7568 34868 7590
rect 2406 7392 2412 7404
rect 2367 7364 2412 7392
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6604 7364 6653 7392
rect 6604 7352 6610 7364
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 20990 7392 20996 7404
rect 20763 7364 20996 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 20990 7352 20996 7364
rect 21048 7352 21054 7404
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 2958 7324 2964 7336
rect 2639 7296 2964 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 6549 7191 6607 7197
rect 6549 7157 6561 7191
rect 6595 7188 6607 7191
rect 7098 7188 7104 7200
rect 6595 7160 7104 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 32674 7188 32680 7200
rect 32635 7160 32680 7188
rect 32674 7148 32680 7160
rect 32732 7148 32738 7200
rect 1104 7098 34868 7120
rect 1104 7046 5174 7098
rect 5226 7046 5238 7098
rect 5290 7046 5302 7098
rect 5354 7046 5366 7098
rect 5418 7046 5430 7098
rect 5482 7046 13622 7098
rect 13674 7046 13686 7098
rect 13738 7046 13750 7098
rect 13802 7046 13814 7098
rect 13866 7046 13878 7098
rect 13930 7046 22070 7098
rect 22122 7046 22134 7098
rect 22186 7046 22198 7098
rect 22250 7046 22262 7098
rect 22314 7046 22326 7098
rect 22378 7046 30518 7098
rect 30570 7046 30582 7098
rect 30634 7046 30646 7098
rect 30698 7046 30710 7098
rect 30762 7046 30774 7098
rect 30826 7046 34868 7098
rect 1104 7024 34868 7046
rect 2958 6848 2964 6860
rect 2919 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7340 6820 8033 6848
rect 7340 6808 7346 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 20070 6848 20076 6860
rect 20031 6820 20076 6848
rect 8021 6811 8079 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 20257 6851 20315 6857
rect 20257 6817 20269 6851
rect 20303 6848 20315 6851
rect 20806 6848 20812 6860
rect 20303 6820 20812 6848
rect 20303 6817 20315 6820
rect 20257 6811 20315 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 21453 6851 21511 6857
rect 21453 6817 21465 6851
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 32309 6851 32367 6857
rect 32309 6817 32321 6851
rect 32355 6848 32367 6851
rect 32674 6848 32680 6860
rect 32355 6820 32680 6848
rect 32355 6817 32367 6820
rect 32309 6811 32367 6817
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10192 6752 10241 6780
rect 10192 6740 10198 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 12802 6780 12808 6792
rect 12763 6752 12808 6780
rect 10229 6743 10287 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13495 6752 14105 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 14093 6749 14105 6752
rect 14139 6780 14151 6783
rect 19702 6780 19708 6792
rect 14139 6752 19708 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 6178 6712 6184 6724
rect 6139 6684 6184 6712
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 7098 6672 7104 6724
rect 7156 6712 7162 6724
rect 7837 6715 7895 6721
rect 7837 6712 7849 6715
rect 7156 6684 7849 6712
rect 7156 6672 7162 6684
rect 7837 6681 7849 6684
rect 7883 6681 7895 6715
rect 7837 6675 7895 6681
rect 20622 6672 20628 6724
rect 20680 6712 20686 6724
rect 21468 6712 21496 6811
rect 32674 6808 32680 6820
rect 32732 6808 32738 6860
rect 34146 6848 34152 6860
rect 34107 6820 34152 6848
rect 34146 6808 34152 6820
rect 34204 6808 34210 6860
rect 27246 6780 27252 6792
rect 27207 6752 27252 6780
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 30561 6783 30619 6789
rect 30561 6749 30573 6783
rect 30607 6780 30619 6783
rect 30926 6780 30932 6792
rect 30607 6752 30932 6780
rect 30607 6749 30619 6752
rect 30561 6743 30619 6749
rect 30926 6740 30932 6752
rect 30984 6740 30990 6792
rect 31202 6780 31208 6792
rect 31163 6752 31208 6780
rect 31202 6740 31208 6752
rect 31260 6740 31266 6792
rect 20680 6684 21496 6712
rect 32493 6715 32551 6721
rect 20680 6672 20686 6684
rect 32493 6681 32505 6715
rect 32539 6712 32551 6715
rect 32582 6712 32588 6724
rect 32539 6684 32588 6712
rect 32539 6681 32551 6684
rect 32493 6675 32551 6681
rect 32582 6672 32588 6684
rect 32640 6672 32646 6724
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 9766 6644 9772 6656
rect 9723 6616 9772 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 12986 6604 12992 6656
rect 13044 6644 13050 6656
rect 13357 6647 13415 6653
rect 13357 6644 13369 6647
rect 13044 6616 13369 6644
rect 13044 6604 13050 6616
rect 13357 6613 13369 6616
rect 13403 6613 13415 6647
rect 13357 6607 13415 6613
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 15746 6644 15752 6656
rect 14231 6616 15752 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 30653 6647 30711 6653
rect 30653 6613 30665 6647
rect 30699 6644 30711 6647
rect 30926 6644 30932 6656
rect 30699 6616 30932 6644
rect 30699 6613 30711 6616
rect 30653 6607 30711 6613
rect 30926 6604 30932 6616
rect 30984 6604 30990 6656
rect 1104 6554 34868 6576
rect 1104 6502 9398 6554
rect 9450 6502 9462 6554
rect 9514 6502 9526 6554
rect 9578 6502 9590 6554
rect 9642 6502 9654 6554
rect 9706 6502 17846 6554
rect 17898 6502 17910 6554
rect 17962 6502 17974 6554
rect 18026 6502 18038 6554
rect 18090 6502 18102 6554
rect 18154 6502 26294 6554
rect 26346 6502 26358 6554
rect 26410 6502 26422 6554
rect 26474 6502 26486 6554
rect 26538 6502 26550 6554
rect 26602 6502 34868 6554
rect 1104 6480 34868 6502
rect 18874 6440 18880 6452
rect 10704 6412 18880 6440
rect 10704 6316 10732 6412
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 32582 6440 32588 6452
rect 32543 6412 32588 6440
rect 32582 6400 32588 6412
rect 32640 6400 32646 6452
rect 12986 6372 12992 6384
rect 12947 6344 12992 6372
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 17126 6332 17132 6384
rect 17184 6372 17190 6384
rect 32122 6372 32128 6384
rect 17184 6344 32128 6372
rect 17184 6332 17190 6344
rect 32122 6332 32128 6344
rect 32180 6372 32186 6384
rect 32398 6372 32404 6384
rect 32180 6344 32404 6372
rect 32180 6332 32186 6344
rect 32398 6332 32404 6344
rect 32456 6332 32462 6384
rect 10686 6304 10692 6316
rect 10599 6276 10692 6304
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 12802 6304 12808 6316
rect 12763 6276 12808 6304
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 27246 6304 27252 6316
rect 27207 6276 27252 6304
rect 27246 6264 27252 6276
rect 27304 6264 27310 6316
rect 32416 6304 32444 6332
rect 32493 6307 32551 6313
rect 32493 6304 32505 6307
rect 32416 6276 32505 6304
rect 32493 6273 32505 6276
rect 32539 6273 32551 6307
rect 32493 6267 32551 6273
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7515 6208 7941 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 8110 6236 8116 6248
rect 8071 6208 8116 6236
rect 7929 6199 7987 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6205 8447 6239
rect 13262 6236 13268 6248
rect 13223 6208 13268 6236
rect 8389 6199 8447 6205
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 8404 6168 8432 6199
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 26970 6196 26976 6248
rect 27028 6236 27034 6248
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 27028 6208 27445 6236
rect 27028 6196 27034 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 29086 6236 29092 6248
rect 29047 6208 29092 6236
rect 27433 6199 27491 6205
rect 29086 6196 29092 6208
rect 29144 6196 29150 6248
rect 5684 6140 8432 6168
rect 5684 6128 5690 6140
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10376 6072 10609 6100
rect 10376 6060 10382 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 15289 6103 15347 6109
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 15930 6100 15936 6112
rect 15335 6072 15936 6100
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 1104 6010 34868 6032
rect 1104 5958 5174 6010
rect 5226 5958 5238 6010
rect 5290 5958 5302 6010
rect 5354 5958 5366 6010
rect 5418 5958 5430 6010
rect 5482 5958 13622 6010
rect 13674 5958 13686 6010
rect 13738 5958 13750 6010
rect 13802 5958 13814 6010
rect 13866 5958 13878 6010
rect 13930 5958 22070 6010
rect 22122 5958 22134 6010
rect 22186 5958 22198 6010
rect 22250 5958 22262 6010
rect 22314 5958 22326 6010
rect 22378 5958 30518 6010
rect 30570 5958 30582 6010
rect 30634 5958 30646 6010
rect 30698 5958 30710 6010
rect 30762 5958 30774 6010
rect 30826 5958 34868 6010
rect 1104 5936 34868 5958
rect 26970 5896 26976 5908
rect 26931 5868 26976 5896
rect 26970 5856 26976 5868
rect 27028 5856 27034 5908
rect 31202 5828 31208 5840
rect 30668 5800 31208 5828
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7098 5760 7104 5772
rect 6595 5732 7104 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 10134 5760 10140 5772
rect 10095 5732 10140 5760
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 10318 5760 10324 5772
rect 10279 5732 10324 5760
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10594 5760 10600 5772
rect 10555 5732 10600 5760
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 15746 5760 15752 5772
rect 15707 5732 15752 5760
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 30668 5769 30696 5800
rect 31202 5788 31208 5800
rect 31260 5788 31266 5840
rect 30653 5763 30711 5769
rect 30653 5729 30665 5763
rect 30699 5729 30711 5763
rect 30653 5723 30711 5729
rect 30837 5763 30895 5769
rect 30837 5729 30849 5763
rect 30883 5760 30895 5763
rect 30926 5760 30932 5772
rect 30883 5732 30932 5760
rect 30883 5729 30895 5732
rect 30837 5723 30895 5729
rect 30926 5720 30932 5732
rect 30984 5720 30990 5772
rect 32214 5760 32220 5772
rect 32175 5732 32220 5760
rect 32214 5720 32220 5732
rect 32272 5720 32278 5772
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 9088 5664 9137 5692
rect 9088 5652 9094 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 19702 5652 19708 5704
rect 19760 5692 19766 5704
rect 26881 5695 26939 5701
rect 26881 5692 26893 5695
rect 19760 5664 26893 5692
rect 19760 5652 19766 5664
rect 26881 5661 26893 5664
rect 26927 5661 26939 5695
rect 27614 5692 27620 5704
rect 27575 5664 27620 5692
rect 26881 5655 26939 5661
rect 27614 5652 27620 5664
rect 27672 5652 27678 5704
rect 6733 5627 6791 5633
rect 6733 5593 6745 5627
rect 6779 5624 6791 5627
rect 7926 5624 7932 5636
rect 6779 5596 7932 5624
rect 6779 5593 6791 5596
rect 6733 5587 6791 5593
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 8386 5624 8392 5636
rect 8347 5596 8392 5624
rect 8386 5584 8392 5596
rect 8444 5584 8450 5636
rect 13538 5584 13544 5636
rect 13596 5624 13602 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 13596 5596 14105 5624
rect 13596 5584 13602 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 14093 5587 14151 5593
rect 1104 5466 34868 5488
rect 1104 5414 9398 5466
rect 9450 5414 9462 5466
rect 9514 5414 9526 5466
rect 9578 5414 9590 5466
rect 9642 5414 9654 5466
rect 9706 5414 17846 5466
rect 17898 5414 17910 5466
rect 17962 5414 17974 5466
rect 18026 5414 18038 5466
rect 18090 5414 18102 5466
rect 18154 5414 26294 5466
rect 26346 5414 26358 5466
rect 26410 5414 26422 5466
rect 26474 5414 26486 5466
rect 26538 5414 26550 5466
rect 26602 5414 34868 5466
rect 1104 5392 34868 5414
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8110 5352 8116 5364
rect 7883 5324 8116 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 10594 5352 10600 5364
rect 9140 5324 10600 5352
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 9140 5284 9168 5324
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 27614 5312 27620 5364
rect 27672 5312 27678 5364
rect 3476 5256 9168 5284
rect 9217 5287 9275 5293
rect 3476 5244 3482 5256
rect 9217 5253 9229 5287
rect 9263 5284 9275 5287
rect 9766 5284 9772 5296
rect 9263 5256 9772 5284
rect 9263 5253 9275 5256
rect 9217 5247 9275 5253
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 27632 5284 27660 5312
rect 27540 5256 27660 5284
rect 7098 5216 7104 5228
rect 7059 5188 7104 5216
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 7929 5179 7987 5185
rect 7944 5148 7972 5179
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 17126 5216 17132 5228
rect 11747 5188 17132 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 27540 5225 27568 5256
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5185 27583 5219
rect 27525 5179 27583 5185
rect 30285 5219 30343 5225
rect 30285 5185 30297 5219
rect 30331 5216 30343 5219
rect 30374 5216 30380 5228
rect 30331 5188 30380 5216
rect 30331 5185 30343 5188
rect 30285 5179 30343 5185
rect 30374 5176 30380 5188
rect 30432 5176 30438 5228
rect 10686 5148 10692 5160
rect 7944 5120 10692 5148
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 10781 5151 10839 5157
rect 10781 5117 10793 5151
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 10796 5080 10824 5111
rect 27338 5108 27344 5160
rect 27396 5148 27402 5160
rect 27709 5151 27767 5157
rect 27709 5148 27721 5151
rect 27396 5120 27721 5148
rect 27396 5108 27402 5120
rect 27709 5117 27721 5120
rect 27755 5117 27767 5151
rect 27709 5111 27767 5117
rect 29365 5151 29423 5157
rect 29365 5117 29377 5151
rect 29411 5148 29423 5151
rect 32306 5148 32312 5160
rect 29411 5120 32312 5148
rect 29411 5117 29423 5120
rect 29365 5111 29423 5117
rect 32306 5108 32312 5120
rect 32364 5108 32370 5160
rect 8260 5052 10824 5080
rect 8260 5040 8266 5052
rect 29086 5040 29092 5092
rect 29144 5080 29150 5092
rect 32398 5080 32404 5092
rect 29144 5052 32404 5080
rect 29144 5040 29150 5052
rect 32398 5040 32404 5052
rect 32456 5040 32462 5092
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7098 5012 7104 5024
rect 6687 4984 7104 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 8573 5015 8631 5021
rect 8573 4981 8585 5015
rect 8619 5012 8631 5015
rect 11146 5012 11152 5024
rect 8619 4984 11152 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11606 5012 11612 5024
rect 11567 4984 11612 5012
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 30374 5012 30380 5024
rect 30335 4984 30380 5012
rect 30374 4972 30380 4984
rect 30432 4972 30438 5024
rect 1104 4922 34868 4944
rect 1104 4870 5174 4922
rect 5226 4870 5238 4922
rect 5290 4870 5302 4922
rect 5354 4870 5366 4922
rect 5418 4870 5430 4922
rect 5482 4870 13622 4922
rect 13674 4870 13686 4922
rect 13738 4870 13750 4922
rect 13802 4870 13814 4922
rect 13866 4870 13878 4922
rect 13930 4870 22070 4922
rect 22122 4870 22134 4922
rect 22186 4870 22198 4922
rect 22250 4870 22262 4922
rect 22314 4870 22326 4922
rect 22378 4870 30518 4922
rect 30570 4870 30582 4922
rect 30634 4870 30646 4922
rect 30698 4870 30710 4922
rect 30762 4870 30774 4922
rect 30826 4870 34868 4922
rect 1104 4848 34868 4870
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 13262 4808 13268 4820
rect 8772 4780 13268 4808
rect 3418 4700 3424 4752
rect 3476 4740 3482 4752
rect 8772 4740 8800 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 27338 4808 27344 4820
rect 27299 4780 27344 4808
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 11606 4740 11612 4752
rect 3476 4712 8800 4740
rect 10980 4712 11612 4740
rect 3476 4700 3482 4712
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 10980 4681 11008 4712
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 30374 4700 30380 4752
rect 30432 4700 30438 4752
rect 10965 4675 11023 4681
rect 6696 4644 8064 4672
rect 6696 4632 6702 4644
rect 7374 4604 7380 4616
rect 7287 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4604 7438 4616
rect 7650 4604 7656 4616
rect 7432 4576 7656 4604
rect 7432 4564 7438 4576
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8036 4613 8064 4644
rect 10965 4641 10977 4675
rect 11011 4641 11023 4675
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 10965 4635 11023 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 30392 4672 30420 4700
rect 30469 4675 30527 4681
rect 30469 4672 30481 4675
rect 30392 4644 30481 4672
rect 30469 4641 30481 4644
rect 30515 4641 30527 4675
rect 30926 4672 30932 4684
rect 30887 4644 30932 4672
rect 30469 4635 30527 4641
rect 30926 4632 30932 4644
rect 30984 4632 30990 4684
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 25314 4564 25320 4616
rect 25372 4604 25378 4616
rect 27249 4607 27307 4613
rect 27249 4604 27261 4607
rect 25372 4576 27261 4604
rect 25372 4564 25378 4576
rect 27249 4573 27261 4576
rect 27295 4573 27307 4607
rect 30282 4604 30288 4616
rect 30243 4576 30288 4604
rect 27249 4567 27307 4573
rect 30282 4564 30288 4576
rect 30340 4564 30346 4616
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 5592 4508 9321 4536
rect 5592 4496 5598 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 1104 4378 34868 4400
rect 1104 4326 9398 4378
rect 9450 4326 9462 4378
rect 9514 4326 9526 4378
rect 9578 4326 9590 4378
rect 9642 4326 9654 4378
rect 9706 4326 17846 4378
rect 17898 4326 17910 4378
rect 17962 4326 17974 4378
rect 18026 4326 18038 4378
rect 18090 4326 18102 4378
rect 18154 4326 26294 4378
rect 26346 4326 26358 4378
rect 26410 4326 26422 4378
rect 26474 4326 26486 4378
rect 26538 4326 26550 4378
rect 26602 4326 34868 4378
rect 1104 4304 34868 4326
rect 7282 4196 7288 4208
rect 7243 4168 7288 4196
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 30282 4128 30288 4140
rect 30243 4100 30288 4128
rect 9861 4091 9919 4097
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 7561 4063 7619 4069
rect 3476 4032 7052 4060
rect 3476 4020 3482 4032
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 7024 3992 7052 4032
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7576 3992 7604 4023
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 9876 4060 9904 4091
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 32122 4088 32128 4140
rect 32180 4128 32186 4140
rect 32217 4131 32275 4137
rect 32217 4128 32229 4131
rect 32180 4100 32229 4128
rect 32180 4088 32186 4100
rect 32217 4097 32229 4100
rect 32263 4097 32275 4131
rect 32217 4091 32275 4097
rect 7708 4032 9904 4060
rect 7708 4020 7714 4032
rect 3936 3964 6914 3992
rect 7024 3964 7604 3992
rect 3936 3952 3942 3964
rect 6886 3924 6914 3964
rect 7834 3924 7840 3936
rect 6886 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 32309 3927 32367 3933
rect 32309 3893 32321 3927
rect 32355 3924 32367 3927
rect 32490 3924 32496 3936
rect 32355 3896 32496 3924
rect 32355 3893 32367 3896
rect 32309 3887 32367 3893
rect 32490 3884 32496 3896
rect 32548 3884 32554 3936
rect 32858 3924 32864 3936
rect 32819 3896 32864 3924
rect 32858 3884 32864 3896
rect 32916 3884 32922 3936
rect 1104 3834 34868 3856
rect 1104 3782 5174 3834
rect 5226 3782 5238 3834
rect 5290 3782 5302 3834
rect 5354 3782 5366 3834
rect 5418 3782 5430 3834
rect 5482 3782 13622 3834
rect 13674 3782 13686 3834
rect 13738 3782 13750 3834
rect 13802 3782 13814 3834
rect 13866 3782 13878 3834
rect 13930 3782 22070 3834
rect 22122 3782 22134 3834
rect 22186 3782 22198 3834
rect 22250 3782 22262 3834
rect 22314 3782 22326 3834
rect 22378 3782 30518 3834
rect 30570 3782 30582 3834
rect 30634 3782 30646 3834
rect 30698 3782 30710 3834
rect 30762 3782 30774 3834
rect 30826 3782 34868 3834
rect 1104 3760 34868 3782
rect 10226 3720 10232 3732
rect 6886 3692 10232 3720
rect 5074 3544 5080 3596
rect 5132 3584 5138 3596
rect 6886 3584 6914 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10502 3652 10508 3664
rect 9784 3624 10508 3652
rect 9784 3593 9812 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 32858 3652 32864 3664
rect 32324 3624 32864 3652
rect 5132 3556 6914 3584
rect 9769 3587 9827 3593
rect 5132 3544 5138 3556
rect 9769 3553 9781 3587
rect 9815 3553 9827 3587
rect 9950 3584 9956 3596
rect 9911 3556 9956 3584
rect 9769 3547 9827 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10318 3584 10324 3596
rect 10279 3556 10324 3584
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 16114 3584 16120 3596
rect 16075 3556 16120 3584
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 32324 3593 32352 3624
rect 32858 3612 32864 3624
rect 32916 3612 32922 3664
rect 32309 3587 32367 3593
rect 32309 3553 32321 3587
rect 32355 3553 32367 3587
rect 32490 3584 32496 3596
rect 32451 3556 32496 3584
rect 32309 3547 32367 3553
rect 32490 3544 32496 3556
rect 32548 3544 32554 3596
rect 2774 3516 2780 3528
rect 2735 3488 2780 3516
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 17644 3488 17877 3516
rect 17644 3476 17650 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 15746 3448 15752 3460
rect 15707 3420 15752 3448
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 34149 3451 34207 3457
rect 34149 3417 34161 3451
rect 34195 3448 34207 3451
rect 34790 3448 34796 3460
rect 34195 3420 34796 3448
rect 34195 3417 34207 3420
rect 34149 3411 34207 3417
rect 34790 3408 34796 3420
rect 34848 3408 34854 3460
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 6178 3380 6184 3392
rect 3292 3352 6184 3380
rect 3292 3340 3298 3352
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 1104 3290 34868 3312
rect 1104 3238 9398 3290
rect 9450 3238 9462 3290
rect 9514 3238 9526 3290
rect 9578 3238 9590 3290
rect 9642 3238 9654 3290
rect 9706 3238 17846 3290
rect 17898 3238 17910 3290
rect 17962 3238 17974 3290
rect 18026 3238 18038 3290
rect 18090 3238 18102 3290
rect 18154 3238 26294 3290
rect 26346 3238 26358 3290
rect 26410 3238 26422 3290
rect 26474 3238 26486 3290
rect 26538 3238 26550 3290
rect 26602 3238 34868 3290
rect 1104 3216 34868 3238
rect 17037 3111 17095 3117
rect 17037 3077 17049 3111
rect 17083 3108 17095 3111
rect 17773 3111 17831 3117
rect 17773 3108 17785 3111
rect 17083 3080 17785 3108
rect 17083 3077 17095 3080
rect 17037 3071 17095 3077
rect 17773 3077 17785 3080
rect 17819 3077 17831 3111
rect 17773 3071 17831 3077
rect 2774 3040 2780 3052
rect 2735 3012 2780 3040
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 15562 3040 15568 3052
rect 15523 3012 15568 3040
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16942 3040 16948 3052
rect 16903 3012 16948 3040
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 2958 2972 2964 2984
rect 2919 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 35434 2972 35440 2984
rect 19475 2944 35440 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3252 2904 3280 2935
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 2648 2876 3280 2904
rect 2648 2864 2654 2876
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 8938 2904 8944 2916
rect 3476 2876 8944 2904
rect 3476 2864 3482 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 5534 2836 5540 2848
rect 4580 2808 5540 2836
rect 4580 2796 4586 2808
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 8202 2836 8208 2848
rect 6512 2808 8208 2836
rect 6512 2796 6518 2808
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 1104 2746 34868 2768
rect 1104 2694 5174 2746
rect 5226 2694 5238 2746
rect 5290 2694 5302 2746
rect 5354 2694 5366 2746
rect 5418 2694 5430 2746
rect 5482 2694 13622 2746
rect 13674 2694 13686 2746
rect 13738 2694 13750 2746
rect 13802 2694 13814 2746
rect 13866 2694 13878 2746
rect 13930 2694 22070 2746
rect 22122 2694 22134 2746
rect 22186 2694 22198 2746
rect 22250 2694 22262 2746
rect 22314 2694 22326 2746
rect 22378 2694 30518 2746
rect 30570 2694 30582 2746
rect 30634 2694 30646 2746
rect 30698 2694 30710 2746
rect 30762 2694 30774 2746
rect 30826 2694 34868 2746
rect 1104 2672 34868 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 3016 2604 3157 2632
rect 3016 2592 3022 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 15746 2632 15752 2644
rect 15707 2604 15752 2632
rect 3145 2595 3203 2601
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 31754 2632 31760 2644
rect 16546 2604 31760 2632
rect 13446 2524 13452 2576
rect 13504 2564 13510 2576
rect 16546 2564 16574 2604
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 13504 2536 16574 2564
rect 13504 2524 13510 2536
rect 3050 2388 3056 2440
rect 3108 2428 3114 2440
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3108 2400 3249 2428
rect 3108 2388 3114 2400
rect 3237 2397 3249 2400
rect 3283 2428 3295 2431
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 3283 2400 15669 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 15657 2397 15669 2400
rect 15703 2428 15715 2431
rect 16942 2428 16948 2440
rect 15703 2400 16948 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 5626 2292 5632 2304
rect 3476 2264 5632 2292
rect 3476 2252 3482 2264
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 1104 2202 34868 2224
rect 1104 2150 9398 2202
rect 9450 2150 9462 2202
rect 9514 2150 9526 2202
rect 9578 2150 9590 2202
rect 9642 2150 9654 2202
rect 9706 2150 17846 2202
rect 17898 2150 17910 2202
rect 17962 2150 17974 2202
rect 18026 2150 18038 2202
rect 18090 2150 18102 2202
rect 18154 2150 26294 2202
rect 26346 2150 26358 2202
rect 26410 2150 26422 2202
rect 26474 2150 26486 2202
rect 26538 2150 26550 2202
rect 26602 2150 34868 2202
rect 1104 2128 34868 2150
<< via1 >>
rect 29736 40060 29788 40112
rect 31760 40060 31812 40112
rect 5174 39686 5226 39738
rect 5238 39686 5290 39738
rect 5302 39686 5354 39738
rect 5366 39686 5418 39738
rect 5430 39686 5482 39738
rect 13622 39686 13674 39738
rect 13686 39686 13738 39738
rect 13750 39686 13802 39738
rect 13814 39686 13866 39738
rect 13878 39686 13930 39738
rect 22070 39686 22122 39738
rect 22134 39686 22186 39738
rect 22198 39686 22250 39738
rect 22262 39686 22314 39738
rect 22326 39686 22378 39738
rect 30518 39686 30570 39738
rect 30582 39686 30634 39738
rect 30646 39686 30698 39738
rect 30710 39686 30762 39738
rect 30774 39686 30826 39738
rect 7840 39423 7892 39432
rect 7840 39389 7849 39423
rect 7849 39389 7883 39423
rect 7883 39389 7892 39423
rect 7840 39380 7892 39389
rect 16120 39423 16172 39432
rect 16120 39389 16129 39423
rect 16129 39389 16163 39423
rect 16163 39389 16172 39423
rect 16120 39380 16172 39389
rect 17040 39423 17092 39432
rect 17040 39389 17049 39423
rect 17049 39389 17083 39423
rect 17083 39389 17092 39423
rect 17040 39380 17092 39389
rect 20996 39423 21048 39432
rect 16948 39312 17000 39364
rect 20996 39389 21005 39423
rect 21005 39389 21039 39423
rect 21039 39389 21048 39423
rect 20996 39380 21048 39389
rect 22376 39380 22428 39432
rect 21088 39312 21140 39364
rect 17132 39287 17184 39296
rect 17132 39253 17141 39287
rect 17141 39253 17175 39287
rect 17175 39253 17184 39287
rect 17132 39244 17184 39253
rect 18052 39244 18104 39296
rect 19248 39244 19300 39296
rect 20812 39244 20864 39296
rect 9398 39142 9450 39194
rect 9462 39142 9514 39194
rect 9526 39142 9578 39194
rect 9590 39142 9642 39194
rect 9654 39142 9706 39194
rect 17846 39142 17898 39194
rect 17910 39142 17962 39194
rect 17974 39142 18026 39194
rect 18038 39142 18090 39194
rect 18102 39142 18154 39194
rect 26294 39142 26346 39194
rect 26358 39142 26410 39194
rect 26422 39142 26474 39194
rect 26486 39142 26538 39194
rect 26550 39142 26602 39194
rect 17132 39015 17184 39024
rect 17132 38981 17141 39015
rect 17141 38981 17175 39015
rect 17175 38981 17184 39015
rect 17132 38972 17184 38981
rect 25136 38972 25188 39024
rect 7840 38947 7892 38956
rect 7840 38913 7849 38947
rect 7849 38913 7883 38947
rect 7883 38913 7892 38947
rect 7840 38904 7892 38913
rect 16948 38947 17000 38956
rect 8024 38879 8076 38888
rect 8024 38845 8033 38879
rect 8033 38845 8067 38879
rect 8067 38845 8076 38879
rect 8024 38836 8076 38845
rect 8392 38879 8444 38888
rect 8392 38845 8401 38879
rect 8401 38845 8435 38879
rect 8435 38845 8444 38879
rect 8392 38836 8444 38845
rect 16948 38913 16957 38947
rect 16957 38913 16991 38947
rect 16991 38913 17000 38947
rect 16948 38904 17000 38913
rect 21088 38947 21140 38956
rect 21088 38913 21097 38947
rect 21097 38913 21131 38947
rect 21131 38913 21140 38947
rect 22376 38947 22428 38956
rect 21088 38904 21140 38913
rect 22376 38913 22385 38947
rect 22385 38913 22419 38947
rect 22419 38913 22428 38947
rect 22376 38904 22428 38913
rect 17408 38879 17460 38888
rect 17408 38845 17417 38879
rect 17417 38845 17451 38879
rect 17451 38845 17460 38879
rect 17408 38836 17460 38845
rect 19340 38879 19392 38888
rect 19340 38845 19349 38879
rect 19349 38845 19383 38879
rect 19383 38845 19392 38879
rect 19340 38836 19392 38845
rect 20904 38879 20956 38888
rect 20904 38845 20913 38879
rect 20913 38845 20947 38879
rect 20947 38845 20956 38879
rect 20904 38836 20956 38845
rect 22560 38879 22612 38888
rect 22560 38845 22569 38879
rect 22569 38845 22603 38879
rect 22603 38845 22612 38879
rect 22560 38836 22612 38845
rect 17040 38768 17092 38820
rect 20260 38768 20312 38820
rect 31760 38768 31812 38820
rect 4896 38700 4948 38752
rect 16580 38700 16632 38752
rect 28448 38700 28500 38752
rect 5174 38598 5226 38650
rect 5238 38598 5290 38650
rect 5302 38598 5354 38650
rect 5366 38598 5418 38650
rect 5430 38598 5482 38650
rect 13622 38598 13674 38650
rect 13686 38598 13738 38650
rect 13750 38598 13802 38650
rect 13814 38598 13866 38650
rect 13878 38598 13930 38650
rect 22070 38598 22122 38650
rect 22134 38598 22186 38650
rect 22198 38598 22250 38650
rect 22262 38598 22314 38650
rect 22326 38598 22378 38650
rect 30518 38598 30570 38650
rect 30582 38598 30634 38650
rect 30646 38598 30698 38650
rect 30710 38598 30762 38650
rect 30774 38598 30826 38650
rect 20 38496 72 38548
rect 1308 38496 1360 38548
rect 8024 38539 8076 38548
rect 8024 38505 8033 38539
rect 8033 38505 8067 38539
rect 8067 38505 8076 38539
rect 8024 38496 8076 38505
rect 22560 38496 22612 38548
rect 4068 38428 4120 38480
rect 4896 38403 4948 38412
rect 4896 38369 4905 38403
rect 4905 38369 4939 38403
rect 4939 38369 4948 38403
rect 4896 38360 4948 38369
rect 9036 38428 9088 38480
rect 19340 38428 19392 38480
rect 19984 38428 20036 38480
rect 16120 38360 16172 38412
rect 16580 38403 16632 38412
rect 16580 38369 16589 38403
rect 16589 38369 16623 38403
rect 16623 38369 16632 38403
rect 16856 38403 16908 38412
rect 16580 38360 16632 38369
rect 16856 38369 16865 38403
rect 16865 38369 16899 38403
rect 16899 38369 16908 38403
rect 16856 38360 16908 38369
rect 20996 38360 21048 38412
rect 6736 38292 6788 38344
rect 23480 38292 23532 38344
rect 28264 38292 28316 38344
rect 30288 38292 30340 38344
rect 32312 38292 32364 38344
rect 5540 38224 5592 38276
rect 20812 38224 20864 38276
rect 16212 38156 16264 38208
rect 16856 38156 16908 38208
rect 28632 38199 28684 38208
rect 28632 38165 28641 38199
rect 28641 38165 28675 38199
rect 28675 38165 28684 38199
rect 28632 38156 28684 38165
rect 9398 38054 9450 38106
rect 9462 38054 9514 38106
rect 9526 38054 9578 38106
rect 9590 38054 9642 38106
rect 9654 38054 9706 38106
rect 17846 38054 17898 38106
rect 17910 38054 17962 38106
rect 17974 38054 18026 38106
rect 18038 38054 18090 38106
rect 18102 38054 18154 38106
rect 26294 38054 26346 38106
rect 26358 38054 26410 38106
rect 26422 38054 26474 38106
rect 26486 38054 26538 38106
rect 26550 38054 26602 38106
rect 5540 37995 5592 38004
rect 5540 37961 5549 37995
rect 5549 37961 5583 37995
rect 5583 37961 5592 37995
rect 5540 37952 5592 37961
rect 20904 37952 20956 38004
rect 20076 37884 20128 37936
rect 34060 37952 34112 38004
rect 28632 37927 28684 37936
rect 28632 37893 28641 37927
rect 28641 37893 28675 37927
rect 28675 37893 28684 37927
rect 28632 37884 28684 37893
rect 34152 37927 34204 37936
rect 34152 37893 34161 37927
rect 34161 37893 34195 37927
rect 34195 37893 34204 37927
rect 34152 37884 34204 37893
rect 6736 37816 6788 37868
rect 7104 37816 7156 37868
rect 10416 37816 10468 37868
rect 28264 37816 28316 37868
rect 28448 37859 28500 37868
rect 28448 37825 28457 37859
rect 28457 37825 28491 37859
rect 28491 37825 28500 37859
rect 28448 37816 28500 37825
rect 32312 37859 32364 37868
rect 32312 37825 32321 37859
rect 32321 37825 32355 37859
rect 32355 37825 32364 37859
rect 32312 37816 32364 37825
rect 29000 37791 29052 37800
rect 29000 37757 29009 37791
rect 29009 37757 29043 37791
rect 29043 37757 29052 37791
rect 29000 37748 29052 37757
rect 32496 37791 32548 37800
rect 32496 37757 32505 37791
rect 32505 37757 32539 37791
rect 32539 37757 32548 37791
rect 32496 37748 32548 37757
rect 8392 37612 8444 37664
rect 22468 37612 22520 37664
rect 5174 37510 5226 37562
rect 5238 37510 5290 37562
rect 5302 37510 5354 37562
rect 5366 37510 5418 37562
rect 5430 37510 5482 37562
rect 13622 37510 13674 37562
rect 13686 37510 13738 37562
rect 13750 37510 13802 37562
rect 13814 37510 13866 37562
rect 13878 37510 13930 37562
rect 22070 37510 22122 37562
rect 22134 37510 22186 37562
rect 22198 37510 22250 37562
rect 22262 37510 22314 37562
rect 22326 37510 22378 37562
rect 30518 37510 30570 37562
rect 30582 37510 30634 37562
rect 30646 37510 30698 37562
rect 30710 37510 30762 37562
rect 30774 37510 30826 37562
rect 32496 37451 32548 37460
rect 32496 37417 32505 37451
rect 32505 37417 32539 37451
rect 32539 37417 32548 37451
rect 32496 37408 32548 37417
rect 664 37204 716 37256
rect 8392 37247 8444 37256
rect 8392 37213 8401 37247
rect 8401 37213 8435 37247
rect 8435 37213 8444 37247
rect 8392 37204 8444 37213
rect 18420 37204 18472 37256
rect 22468 37272 22520 37324
rect 22652 37315 22704 37324
rect 22652 37281 22661 37315
rect 22661 37281 22695 37315
rect 22695 37281 22704 37315
rect 22652 37272 22704 37281
rect 30288 37272 30340 37324
rect 7380 37136 7432 37188
rect 22192 37179 22244 37188
rect 22192 37145 22201 37179
rect 22201 37145 22235 37179
rect 22235 37145 22244 37179
rect 22192 37136 22244 37145
rect 9398 36966 9450 37018
rect 9462 36966 9514 37018
rect 9526 36966 9578 37018
rect 9590 36966 9642 37018
rect 9654 36966 9706 37018
rect 17846 36966 17898 37018
rect 17910 36966 17962 37018
rect 17974 36966 18026 37018
rect 18038 36966 18090 37018
rect 18102 36966 18154 37018
rect 26294 36966 26346 37018
rect 26358 36966 26410 37018
rect 26422 36966 26474 37018
rect 26486 36966 26538 37018
rect 26550 36966 26602 37018
rect 7380 36907 7432 36916
rect 7380 36873 7389 36907
rect 7389 36873 7423 36907
rect 7423 36873 7432 36907
rect 7380 36864 7432 36873
rect 22192 36907 22244 36916
rect 22192 36873 22201 36907
rect 22201 36873 22235 36907
rect 22235 36873 22244 36907
rect 22192 36864 22244 36873
rect 20260 36839 20312 36848
rect 20260 36805 20269 36839
rect 20269 36805 20303 36839
rect 20303 36805 20312 36839
rect 20260 36796 20312 36805
rect 17500 36728 17552 36780
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 27804 36728 27856 36780
rect 17316 36567 17368 36576
rect 17316 36533 17325 36567
rect 17325 36533 17359 36567
rect 17359 36533 17368 36567
rect 17316 36524 17368 36533
rect 5174 36422 5226 36474
rect 5238 36422 5290 36474
rect 5302 36422 5354 36474
rect 5366 36422 5418 36474
rect 5430 36422 5482 36474
rect 13622 36422 13674 36474
rect 13686 36422 13738 36474
rect 13750 36422 13802 36474
rect 13814 36422 13866 36474
rect 13878 36422 13930 36474
rect 22070 36422 22122 36474
rect 22134 36422 22186 36474
rect 22198 36422 22250 36474
rect 22262 36422 22314 36474
rect 22326 36422 22378 36474
rect 30518 36422 30570 36474
rect 30582 36422 30634 36474
rect 30646 36422 30698 36474
rect 30710 36422 30762 36474
rect 30774 36422 30826 36474
rect 17500 36159 17552 36168
rect 17500 36125 17509 36159
rect 17509 36125 17543 36159
rect 17543 36125 17552 36159
rect 17500 36116 17552 36125
rect 27896 36159 27948 36168
rect 27896 36125 27905 36159
rect 27905 36125 27939 36159
rect 27939 36125 27948 36159
rect 27896 36116 27948 36125
rect 1860 36091 1912 36100
rect 1860 36057 1869 36091
rect 1869 36057 1903 36091
rect 1903 36057 1912 36091
rect 1860 36048 1912 36057
rect 1952 36023 2004 36032
rect 1952 35989 1961 36023
rect 1961 35989 1995 36023
rect 1995 35989 2004 36023
rect 1952 35980 2004 35989
rect 17684 35980 17736 36032
rect 9398 35878 9450 35930
rect 9462 35878 9514 35930
rect 9526 35878 9578 35930
rect 9590 35878 9642 35930
rect 9654 35878 9706 35930
rect 17846 35878 17898 35930
rect 17910 35878 17962 35930
rect 17974 35878 18026 35930
rect 18038 35878 18090 35930
rect 18102 35878 18154 35930
rect 26294 35878 26346 35930
rect 26358 35878 26410 35930
rect 26422 35878 26474 35930
rect 26486 35878 26538 35930
rect 26550 35878 26602 35930
rect 17684 35751 17736 35760
rect 17684 35717 17693 35751
rect 17693 35717 17727 35751
rect 17727 35717 17736 35751
rect 17684 35708 17736 35717
rect 29736 35751 29788 35760
rect 29736 35717 29745 35751
rect 29745 35717 29779 35751
rect 29779 35717 29788 35751
rect 29736 35708 29788 35717
rect 17316 35640 17368 35692
rect 27896 35683 27948 35692
rect 27896 35649 27905 35683
rect 27905 35649 27939 35683
rect 27939 35649 27948 35683
rect 27896 35640 27948 35649
rect 19248 35615 19300 35624
rect 19248 35581 19257 35615
rect 19257 35581 19291 35615
rect 19291 35581 19300 35615
rect 19248 35572 19300 35581
rect 28080 35615 28132 35624
rect 28080 35581 28089 35615
rect 28089 35581 28123 35615
rect 28123 35581 28132 35615
rect 28080 35572 28132 35581
rect 5174 35334 5226 35386
rect 5238 35334 5290 35386
rect 5302 35334 5354 35386
rect 5366 35334 5418 35386
rect 5430 35334 5482 35386
rect 13622 35334 13674 35386
rect 13686 35334 13738 35386
rect 13750 35334 13802 35386
rect 13814 35334 13866 35386
rect 13878 35334 13930 35386
rect 22070 35334 22122 35386
rect 22134 35334 22186 35386
rect 22198 35334 22250 35386
rect 22262 35334 22314 35386
rect 22326 35334 22378 35386
rect 30518 35334 30570 35386
rect 30582 35334 30634 35386
rect 30646 35334 30698 35386
rect 30710 35334 30762 35386
rect 30774 35334 30826 35386
rect 28080 35232 28132 35284
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 29092 35028 29144 35080
rect 9398 34790 9450 34842
rect 9462 34790 9514 34842
rect 9526 34790 9578 34842
rect 9590 34790 9642 34842
rect 9654 34790 9706 34842
rect 17846 34790 17898 34842
rect 17910 34790 17962 34842
rect 17974 34790 18026 34842
rect 18038 34790 18090 34842
rect 18102 34790 18154 34842
rect 26294 34790 26346 34842
rect 26358 34790 26410 34842
rect 26422 34790 26474 34842
rect 26486 34790 26538 34842
rect 26550 34790 26602 34842
rect 9864 34348 9916 34400
rect 5174 34246 5226 34298
rect 5238 34246 5290 34298
rect 5302 34246 5354 34298
rect 5366 34246 5418 34298
rect 5430 34246 5482 34298
rect 13622 34246 13674 34298
rect 13686 34246 13738 34298
rect 13750 34246 13802 34298
rect 13814 34246 13866 34298
rect 13878 34246 13930 34298
rect 22070 34246 22122 34298
rect 22134 34246 22186 34298
rect 22198 34246 22250 34298
rect 22262 34246 22314 34298
rect 22326 34246 22378 34298
rect 30518 34246 30570 34298
rect 30582 34246 30634 34298
rect 30646 34246 30698 34298
rect 30710 34246 30762 34298
rect 30774 34246 30826 34298
rect 3424 33872 3476 33924
rect 9864 34051 9916 34060
rect 9864 34017 9873 34051
rect 9873 34017 9907 34051
rect 9907 34017 9916 34051
rect 9864 34008 9916 34017
rect 27620 33983 27672 33992
rect 27620 33949 27629 33983
rect 27629 33949 27663 33983
rect 27663 33949 27672 33983
rect 27620 33940 27672 33949
rect 10232 33872 10284 33924
rect 9398 33702 9450 33754
rect 9462 33702 9514 33754
rect 9526 33702 9578 33754
rect 9590 33702 9642 33754
rect 9654 33702 9706 33754
rect 17846 33702 17898 33754
rect 17910 33702 17962 33754
rect 17974 33702 18026 33754
rect 18038 33702 18090 33754
rect 18102 33702 18154 33754
rect 26294 33702 26346 33754
rect 26358 33702 26410 33754
rect 26422 33702 26474 33754
rect 26486 33702 26538 33754
rect 26550 33702 26602 33754
rect 10232 33643 10284 33652
rect 10232 33609 10241 33643
rect 10241 33609 10275 33643
rect 10275 33609 10284 33643
rect 10232 33600 10284 33609
rect 10324 33507 10376 33516
rect 10324 33473 10333 33507
rect 10333 33473 10367 33507
rect 10367 33473 10376 33507
rect 10324 33464 10376 33473
rect 27620 33507 27672 33516
rect 27620 33473 27629 33507
rect 27629 33473 27663 33507
rect 27663 33473 27672 33507
rect 27620 33464 27672 33473
rect 27804 33439 27856 33448
rect 27804 33405 27813 33439
rect 27813 33405 27847 33439
rect 27847 33405 27856 33439
rect 27804 33396 27856 33405
rect 32312 33396 32364 33448
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 5174 33158 5226 33210
rect 5238 33158 5290 33210
rect 5302 33158 5354 33210
rect 5366 33158 5418 33210
rect 5430 33158 5482 33210
rect 13622 33158 13674 33210
rect 13686 33158 13738 33210
rect 13750 33158 13802 33210
rect 13814 33158 13866 33210
rect 13878 33158 13930 33210
rect 22070 33158 22122 33210
rect 22134 33158 22186 33210
rect 22198 33158 22250 33210
rect 22262 33158 22314 33210
rect 22326 33158 22378 33210
rect 30518 33158 30570 33210
rect 30582 33158 30634 33210
rect 30646 33158 30698 33210
rect 30710 33158 30762 33210
rect 30774 33158 30826 33210
rect 27804 33056 27856 33108
rect 17040 32920 17092 32972
rect 18236 32852 18288 32904
rect 32128 32920 32180 32972
rect 29828 32852 29880 32904
rect 30288 32852 30340 32904
rect 33692 32827 33744 32836
rect 33692 32793 33701 32827
rect 33701 32793 33735 32827
rect 33735 32793 33744 32827
rect 33692 32784 33744 32793
rect 9398 32614 9450 32666
rect 9462 32614 9514 32666
rect 9526 32614 9578 32666
rect 9590 32614 9642 32666
rect 9654 32614 9706 32666
rect 17846 32614 17898 32666
rect 17910 32614 17962 32666
rect 17974 32614 18026 32666
rect 18038 32614 18090 32666
rect 18102 32614 18154 32666
rect 26294 32614 26346 32666
rect 26358 32614 26410 32666
rect 26422 32614 26474 32666
rect 26486 32614 26538 32666
rect 26550 32614 26602 32666
rect 20076 32487 20128 32496
rect 20076 32453 20085 32487
rect 20085 32453 20119 32487
rect 20119 32453 20128 32487
rect 20076 32444 20128 32453
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 17960 32308 18012 32360
rect 32312 32351 32364 32360
rect 32312 32317 32321 32351
rect 32321 32317 32355 32351
rect 32355 32317 32364 32351
rect 32312 32308 32364 32317
rect 31852 32240 31904 32292
rect 5174 32070 5226 32122
rect 5238 32070 5290 32122
rect 5302 32070 5354 32122
rect 5366 32070 5418 32122
rect 5430 32070 5482 32122
rect 13622 32070 13674 32122
rect 13686 32070 13738 32122
rect 13750 32070 13802 32122
rect 13814 32070 13866 32122
rect 13878 32070 13930 32122
rect 22070 32070 22122 32122
rect 22134 32070 22186 32122
rect 22198 32070 22250 32122
rect 22262 32070 22314 32122
rect 22326 32070 22378 32122
rect 30518 32070 30570 32122
rect 30582 32070 30634 32122
rect 30646 32070 30698 32122
rect 30710 32070 30762 32122
rect 30774 32070 30826 32122
rect 17960 32011 18012 32020
rect 17960 31977 17969 32011
rect 17969 31977 18003 32011
rect 18003 31977 18012 32011
rect 17960 31968 18012 31977
rect 32312 31968 32364 32020
rect 17040 31832 17092 31884
rect 17592 31832 17644 31884
rect 19524 31832 19576 31884
rect 3424 31764 3476 31816
rect 10968 31764 11020 31816
rect 16304 31764 16356 31816
rect 26976 31764 27028 31816
rect 32036 31764 32088 31816
rect 20260 31739 20312 31748
rect 20260 31705 20269 31739
rect 20269 31705 20303 31739
rect 20303 31705 20312 31739
rect 20260 31696 20312 31705
rect 9398 31526 9450 31578
rect 9462 31526 9514 31578
rect 9526 31526 9578 31578
rect 9590 31526 9642 31578
rect 9654 31526 9706 31578
rect 17846 31526 17898 31578
rect 17910 31526 17962 31578
rect 17974 31526 18026 31578
rect 18038 31526 18090 31578
rect 18102 31526 18154 31578
rect 26294 31526 26346 31578
rect 26358 31526 26410 31578
rect 26422 31526 26474 31578
rect 26486 31526 26538 31578
rect 26550 31526 26602 31578
rect 20260 31467 20312 31476
rect 20260 31433 20269 31467
rect 20269 31433 20303 31467
rect 20303 31433 20312 31467
rect 20260 31424 20312 31433
rect 20168 31331 20220 31340
rect 20168 31297 20177 31331
rect 20177 31297 20211 31331
rect 20211 31297 20220 31331
rect 20168 31288 20220 31297
rect 24860 31288 24912 31340
rect 26976 31331 27028 31340
rect 26976 31297 26985 31331
rect 26985 31297 27019 31331
rect 27019 31297 27028 31331
rect 26976 31288 27028 31297
rect 20 31220 72 31272
rect 11704 31263 11756 31272
rect 11704 31229 11713 31263
rect 11713 31229 11747 31263
rect 11747 31229 11756 31263
rect 11704 31220 11756 31229
rect 26700 31152 26752 31204
rect 5174 30982 5226 31034
rect 5238 30982 5290 31034
rect 5302 30982 5354 31034
rect 5366 30982 5418 31034
rect 5430 30982 5482 31034
rect 13622 30982 13674 31034
rect 13686 30982 13738 31034
rect 13750 30982 13802 31034
rect 13814 30982 13866 31034
rect 13878 30982 13930 31034
rect 22070 30982 22122 31034
rect 22134 30982 22186 31034
rect 22198 30982 22250 31034
rect 22262 30982 22314 31034
rect 22326 30982 22378 31034
rect 30518 30982 30570 31034
rect 30582 30982 30634 31034
rect 30646 30982 30698 31034
rect 30710 30982 30762 31034
rect 30774 30982 30826 31034
rect 11704 30880 11756 30932
rect 2780 30676 2832 30728
rect 11796 30676 11848 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 33968 30719 34020 30728
rect 33968 30685 33977 30719
rect 33977 30685 34011 30719
rect 34011 30685 34020 30719
rect 33968 30676 34020 30685
rect 18236 30608 18288 30660
rect 9398 30438 9450 30490
rect 9462 30438 9514 30490
rect 9526 30438 9578 30490
rect 9590 30438 9642 30490
rect 9654 30438 9706 30490
rect 17846 30438 17898 30490
rect 17910 30438 17962 30490
rect 17974 30438 18026 30490
rect 18038 30438 18090 30490
rect 18102 30438 18154 30490
rect 26294 30438 26346 30490
rect 26358 30438 26410 30490
rect 26422 30438 26474 30490
rect 26486 30438 26538 30490
rect 26550 30438 26602 30490
rect 20168 30336 20220 30388
rect 27804 30336 27856 30388
rect 2780 30243 2832 30252
rect 2780 30209 2789 30243
rect 2789 30209 2823 30243
rect 2823 30209 2832 30243
rect 2780 30200 2832 30209
rect 11796 30243 11848 30252
rect 11796 30209 11805 30243
rect 11805 30209 11839 30243
rect 11839 30209 11848 30243
rect 11796 30200 11848 30209
rect 14280 30243 14332 30252
rect 14280 30209 14289 30243
rect 14289 30209 14323 30243
rect 14323 30209 14332 30243
rect 14280 30200 14332 30209
rect 3148 30132 3200 30184
rect 4160 30175 4212 30184
rect 4160 30141 4169 30175
rect 4169 30141 4203 30175
rect 4203 30141 4212 30175
rect 4160 30132 4212 30141
rect 12164 30132 12216 30184
rect 14464 30175 14516 30184
rect 10968 30064 11020 30116
rect 14464 30141 14473 30175
rect 14473 30141 14507 30175
rect 14507 30141 14516 30175
rect 14464 30132 14516 30141
rect 14832 30175 14884 30184
rect 14832 30141 14841 30175
rect 14841 30141 14875 30175
rect 14875 30141 14884 30175
rect 14832 30132 14884 30141
rect 19340 29996 19392 30048
rect 27068 29996 27120 30048
rect 32312 29996 32364 30048
rect 33784 30039 33836 30048
rect 33784 30005 33793 30039
rect 33793 30005 33827 30039
rect 33827 30005 33836 30039
rect 33784 29996 33836 30005
rect 5174 29894 5226 29946
rect 5238 29894 5290 29946
rect 5302 29894 5354 29946
rect 5366 29894 5418 29946
rect 5430 29894 5482 29946
rect 13622 29894 13674 29946
rect 13686 29894 13738 29946
rect 13750 29894 13802 29946
rect 13814 29894 13866 29946
rect 13878 29894 13930 29946
rect 22070 29894 22122 29946
rect 22134 29894 22186 29946
rect 22198 29894 22250 29946
rect 22262 29894 22314 29946
rect 22326 29894 22378 29946
rect 30518 29894 30570 29946
rect 30582 29894 30634 29946
rect 30646 29894 30698 29946
rect 30710 29894 30762 29946
rect 30774 29894 30826 29946
rect 3148 29835 3200 29844
rect 3148 29801 3157 29835
rect 3157 29801 3191 29835
rect 3191 29801 3200 29835
rect 3148 29792 3200 29801
rect 12164 29835 12216 29844
rect 12164 29801 12173 29835
rect 12173 29801 12207 29835
rect 12207 29801 12216 29835
rect 12164 29792 12216 29801
rect 14464 29835 14516 29844
rect 14464 29801 14473 29835
rect 14473 29801 14507 29835
rect 14507 29801 14516 29835
rect 14464 29792 14516 29801
rect 2964 29588 3016 29640
rect 3424 29520 3476 29572
rect 19340 29699 19392 29708
rect 19340 29665 19349 29699
rect 19349 29665 19383 29699
rect 19383 29665 19392 29699
rect 19340 29656 19392 29665
rect 25412 29656 25464 29708
rect 33048 29699 33100 29708
rect 33048 29665 33057 29699
rect 33057 29665 33091 29699
rect 33091 29665 33100 29699
rect 33048 29656 33100 29665
rect 33968 29656 34020 29708
rect 16304 29588 16356 29640
rect 25228 29631 25280 29640
rect 25228 29597 25237 29631
rect 25237 29597 25271 29631
rect 25271 29597 25280 29631
rect 25228 29588 25280 29597
rect 19800 29520 19852 29572
rect 25412 29563 25464 29572
rect 25412 29529 25421 29563
rect 25421 29529 25455 29563
rect 25455 29529 25464 29563
rect 25412 29520 25464 29529
rect 29368 29588 29420 29640
rect 33968 29563 34020 29572
rect 19340 29452 19392 29504
rect 20720 29452 20772 29504
rect 33968 29529 33977 29563
rect 33977 29529 34011 29563
rect 34011 29529 34020 29563
rect 33968 29520 34020 29529
rect 27252 29452 27304 29504
rect 9398 29350 9450 29402
rect 9462 29350 9514 29402
rect 9526 29350 9578 29402
rect 9590 29350 9642 29402
rect 9654 29350 9706 29402
rect 17846 29350 17898 29402
rect 17910 29350 17962 29402
rect 17974 29350 18026 29402
rect 18038 29350 18090 29402
rect 18102 29350 18154 29402
rect 26294 29350 26346 29402
rect 26358 29350 26410 29402
rect 26422 29350 26474 29402
rect 26486 29350 26538 29402
rect 26550 29350 26602 29402
rect 2964 29248 3016 29300
rect 18328 29248 18380 29300
rect 19800 29291 19852 29300
rect 19800 29257 19809 29291
rect 19809 29257 19843 29291
rect 19843 29257 19852 29291
rect 19800 29248 19852 29257
rect 27252 29223 27304 29232
rect 27252 29189 27261 29223
rect 27261 29189 27295 29223
rect 27295 29189 27304 29223
rect 27252 29180 27304 29189
rect 31668 29180 31720 29232
rect 34152 29223 34204 29232
rect 34152 29189 34161 29223
rect 34161 29189 34195 29223
rect 34195 29189 34204 29223
rect 34152 29180 34204 29189
rect 20720 29112 20772 29164
rect 25228 29112 25280 29164
rect 27068 29155 27120 29164
rect 27068 29121 27077 29155
rect 27077 29121 27111 29155
rect 27111 29121 27120 29155
rect 27068 29112 27120 29121
rect 29368 29155 29420 29164
rect 29368 29121 29377 29155
rect 29377 29121 29411 29155
rect 29411 29121 29420 29155
rect 29368 29112 29420 29121
rect 32312 29155 32364 29164
rect 32312 29121 32321 29155
rect 32321 29121 32355 29155
rect 32355 29121 32364 29155
rect 32312 29112 32364 29121
rect 28448 29087 28500 29096
rect 28448 29053 28457 29087
rect 28457 29053 28491 29087
rect 28491 29053 28500 29087
rect 28448 29044 28500 29053
rect 29552 29087 29604 29096
rect 29552 29053 29561 29087
rect 29561 29053 29595 29087
rect 29595 29053 29604 29087
rect 29552 29044 29604 29053
rect 32496 29087 32548 29096
rect 32496 29053 32505 29087
rect 32505 29053 32539 29087
rect 32539 29053 32548 29087
rect 32496 29044 32548 29053
rect 25504 28951 25556 28960
rect 25504 28917 25513 28951
rect 25513 28917 25547 28951
rect 25547 28917 25556 28951
rect 25504 28908 25556 28917
rect 5174 28806 5226 28858
rect 5238 28806 5290 28858
rect 5302 28806 5354 28858
rect 5366 28806 5418 28858
rect 5430 28806 5482 28858
rect 13622 28806 13674 28858
rect 13686 28806 13738 28858
rect 13750 28806 13802 28858
rect 13814 28806 13866 28858
rect 13878 28806 13930 28858
rect 22070 28806 22122 28858
rect 22134 28806 22186 28858
rect 22198 28806 22250 28858
rect 22262 28806 22314 28858
rect 22326 28806 22378 28858
rect 30518 28806 30570 28858
rect 30582 28806 30634 28858
rect 30646 28806 30698 28858
rect 30710 28806 30762 28858
rect 30774 28806 30826 28858
rect 25412 28704 25464 28756
rect 29552 28704 29604 28756
rect 25504 28611 25556 28620
rect 25504 28577 25513 28611
rect 25513 28577 25547 28611
rect 25547 28577 25556 28611
rect 25504 28568 25556 28577
rect 31576 28568 31628 28620
rect 33508 28611 33560 28620
rect 33508 28577 33517 28611
rect 33517 28577 33551 28611
rect 33551 28577 33560 28611
rect 33508 28568 33560 28577
rect 33784 28568 33836 28620
rect 19708 28500 19760 28552
rect 24860 28543 24912 28552
rect 24860 28509 24869 28543
rect 24869 28509 24903 28543
rect 24903 28509 24912 28543
rect 24860 28500 24912 28509
rect 27804 28543 27856 28552
rect 27804 28509 27813 28543
rect 27813 28509 27847 28543
rect 27847 28509 27856 28543
rect 27804 28500 27856 28509
rect 25504 28432 25556 28484
rect 33416 28432 33468 28484
rect 9398 28262 9450 28314
rect 9462 28262 9514 28314
rect 9526 28262 9578 28314
rect 9590 28262 9642 28314
rect 9654 28262 9706 28314
rect 17846 28262 17898 28314
rect 17910 28262 17962 28314
rect 17974 28262 18026 28314
rect 18038 28262 18090 28314
rect 18102 28262 18154 28314
rect 26294 28262 26346 28314
rect 26358 28262 26410 28314
rect 26422 28262 26474 28314
rect 26486 28262 26538 28314
rect 26550 28262 26602 28314
rect 25504 28203 25556 28212
rect 25504 28169 25513 28203
rect 25513 28169 25547 28203
rect 25547 28169 25556 28203
rect 25504 28160 25556 28169
rect 32496 28160 32548 28212
rect 33416 28203 33468 28212
rect 33416 28169 33425 28203
rect 33425 28169 33459 28203
rect 33459 28169 33468 28203
rect 33416 28160 33468 28169
rect 33968 28160 34020 28212
rect 25412 28067 25464 28076
rect 25412 28033 25421 28067
rect 25421 28033 25455 28067
rect 25455 28033 25464 28067
rect 25412 28024 25464 28033
rect 33140 28024 33192 28076
rect 33324 28024 33376 28076
rect 5174 27718 5226 27770
rect 5238 27718 5290 27770
rect 5302 27718 5354 27770
rect 5366 27718 5418 27770
rect 5430 27718 5482 27770
rect 13622 27718 13674 27770
rect 13686 27718 13738 27770
rect 13750 27718 13802 27770
rect 13814 27718 13866 27770
rect 13878 27718 13930 27770
rect 22070 27718 22122 27770
rect 22134 27718 22186 27770
rect 22198 27718 22250 27770
rect 22262 27718 22314 27770
rect 22326 27718 22378 27770
rect 30518 27718 30570 27770
rect 30582 27718 30634 27770
rect 30646 27718 30698 27770
rect 30710 27718 30762 27770
rect 30774 27718 30826 27770
rect 9398 27174 9450 27226
rect 9462 27174 9514 27226
rect 9526 27174 9578 27226
rect 9590 27174 9642 27226
rect 9654 27174 9706 27226
rect 17846 27174 17898 27226
rect 17910 27174 17962 27226
rect 17974 27174 18026 27226
rect 18038 27174 18090 27226
rect 18102 27174 18154 27226
rect 26294 27174 26346 27226
rect 26358 27174 26410 27226
rect 26422 27174 26474 27226
rect 26486 27174 26538 27226
rect 26550 27174 26602 27226
rect 31300 26775 31352 26784
rect 31300 26741 31309 26775
rect 31309 26741 31343 26775
rect 31343 26741 31352 26775
rect 31300 26732 31352 26741
rect 5174 26630 5226 26682
rect 5238 26630 5290 26682
rect 5302 26630 5354 26682
rect 5366 26630 5418 26682
rect 5430 26630 5482 26682
rect 13622 26630 13674 26682
rect 13686 26630 13738 26682
rect 13750 26630 13802 26682
rect 13814 26630 13866 26682
rect 13878 26630 13930 26682
rect 22070 26630 22122 26682
rect 22134 26630 22186 26682
rect 22198 26630 22250 26682
rect 22262 26630 22314 26682
rect 22326 26630 22378 26682
rect 30518 26630 30570 26682
rect 30582 26630 30634 26682
rect 30646 26630 30698 26682
rect 30710 26630 30762 26682
rect 30774 26630 30826 26682
rect 31300 26435 31352 26444
rect 31300 26401 31309 26435
rect 31309 26401 31343 26435
rect 31343 26401 31352 26435
rect 31300 26392 31352 26401
rect 33048 26435 33100 26444
rect 33048 26401 33057 26435
rect 33057 26401 33091 26435
rect 33091 26401 33100 26435
rect 33048 26392 33100 26401
rect 8852 26324 8904 26376
rect 29736 26324 29788 26376
rect 32220 26256 32272 26308
rect 9398 26086 9450 26138
rect 9462 26086 9514 26138
rect 9526 26086 9578 26138
rect 9590 26086 9642 26138
rect 9654 26086 9706 26138
rect 17846 26086 17898 26138
rect 17910 26086 17962 26138
rect 17974 26086 18026 26138
rect 18038 26086 18090 26138
rect 18102 26086 18154 26138
rect 26294 26086 26346 26138
rect 26358 26086 26410 26138
rect 26422 26086 26474 26138
rect 26486 26086 26538 26138
rect 26550 26086 26602 26138
rect 32220 26027 32272 26036
rect 32220 25993 32229 26027
rect 32229 25993 32263 26027
rect 32263 25993 32272 26027
rect 32220 25984 32272 25993
rect 3608 25916 3660 25968
rect 8852 25916 8904 25968
rect 33048 25916 33100 25968
rect 29092 25891 29144 25900
rect 29092 25857 29101 25891
rect 29101 25857 29135 25891
rect 29135 25857 29144 25891
rect 29092 25848 29144 25857
rect 29736 25891 29788 25900
rect 29736 25857 29745 25891
rect 29745 25857 29779 25891
rect 29779 25857 29788 25891
rect 29736 25848 29788 25857
rect 31944 25848 31996 25900
rect 9036 25780 9088 25832
rect 9956 25644 10008 25696
rect 5174 25542 5226 25594
rect 5238 25542 5290 25594
rect 5302 25542 5354 25594
rect 5366 25542 5418 25594
rect 5430 25542 5482 25594
rect 13622 25542 13674 25594
rect 13686 25542 13738 25594
rect 13750 25542 13802 25594
rect 13814 25542 13866 25594
rect 13878 25542 13930 25594
rect 22070 25542 22122 25594
rect 22134 25542 22186 25594
rect 22198 25542 22250 25594
rect 22262 25542 22314 25594
rect 22326 25542 22378 25594
rect 30518 25542 30570 25594
rect 30582 25542 30634 25594
rect 30646 25542 30698 25594
rect 30710 25542 30762 25594
rect 30774 25542 30826 25594
rect 9036 25483 9088 25492
rect 9036 25449 9045 25483
rect 9045 25449 9079 25483
rect 9079 25449 9088 25483
rect 9036 25440 9088 25449
rect 9956 25347 10008 25356
rect 9956 25313 9965 25347
rect 9965 25313 9999 25347
rect 9999 25313 10008 25347
rect 9956 25304 10008 25313
rect 10416 25347 10468 25356
rect 10416 25313 10425 25347
rect 10425 25313 10459 25347
rect 10459 25313 10468 25347
rect 10416 25304 10468 25313
rect 32956 25347 33008 25356
rect 32956 25313 32965 25347
rect 32965 25313 32999 25347
rect 32999 25313 33008 25347
rect 32956 25304 33008 25313
rect 7656 25236 7708 25288
rect 9312 25236 9364 25288
rect 10140 25211 10192 25220
rect 10140 25177 10149 25211
rect 10149 25177 10183 25211
rect 10183 25177 10192 25211
rect 10140 25168 10192 25177
rect 31668 25211 31720 25220
rect 31668 25177 31677 25211
rect 31677 25177 31711 25211
rect 31711 25177 31720 25211
rect 31668 25168 31720 25177
rect 9398 24998 9450 25050
rect 9462 24998 9514 25050
rect 9526 24998 9578 25050
rect 9590 24998 9642 25050
rect 9654 24998 9706 25050
rect 17846 24998 17898 25050
rect 17910 24998 17962 25050
rect 17974 24998 18026 25050
rect 18038 24998 18090 25050
rect 18102 24998 18154 25050
rect 26294 24998 26346 25050
rect 26358 24998 26410 25050
rect 26422 24998 26474 25050
rect 26486 24998 26538 25050
rect 26550 24998 26602 25050
rect 3424 24896 3476 24948
rect 8392 24896 8444 24948
rect 10140 24896 10192 24948
rect 31668 24896 31720 24948
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 11060 24760 11112 24812
rect 18328 24760 18380 24812
rect 25412 24760 25464 24812
rect 27068 24760 27120 24812
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 8300 24692 8352 24744
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 32312 24556 32364 24608
rect 5174 24454 5226 24506
rect 5238 24454 5290 24506
rect 5302 24454 5354 24506
rect 5366 24454 5418 24506
rect 5430 24454 5482 24506
rect 13622 24454 13674 24506
rect 13686 24454 13738 24506
rect 13750 24454 13802 24506
rect 13814 24454 13866 24506
rect 13878 24454 13930 24506
rect 22070 24454 22122 24506
rect 22134 24454 22186 24506
rect 22198 24454 22250 24506
rect 22262 24454 22314 24506
rect 22326 24454 22378 24506
rect 30518 24454 30570 24506
rect 30582 24454 30634 24506
rect 30646 24454 30698 24506
rect 30710 24454 30762 24506
rect 30774 24454 30826 24506
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 11060 24148 11112 24200
rect 29828 24191 29880 24200
rect 19616 24080 19668 24132
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 30932 24148 30984 24200
rect 32036 24148 32088 24200
rect 32772 24191 32824 24200
rect 32772 24157 32781 24191
rect 32781 24157 32815 24191
rect 32815 24157 32824 24191
rect 32772 24148 32824 24157
rect 29920 24055 29972 24064
rect 29920 24021 29929 24055
rect 29929 24021 29963 24055
rect 29963 24021 29972 24055
rect 29920 24012 29972 24021
rect 32496 24012 32548 24064
rect 9398 23910 9450 23962
rect 9462 23910 9514 23962
rect 9526 23910 9578 23962
rect 9590 23910 9642 23962
rect 9654 23910 9706 23962
rect 17846 23910 17898 23962
rect 17910 23910 17962 23962
rect 17974 23910 18026 23962
rect 18038 23910 18090 23962
rect 18102 23910 18154 23962
rect 26294 23910 26346 23962
rect 26358 23910 26410 23962
rect 26422 23910 26474 23962
rect 26486 23910 26538 23962
rect 26550 23910 26602 23962
rect 1952 23672 2004 23724
rect 16580 23672 16632 23724
rect 18328 23740 18380 23792
rect 29920 23783 29972 23792
rect 29920 23749 29929 23783
rect 29929 23749 29963 23783
rect 29963 23749 29972 23783
rect 29920 23740 29972 23749
rect 32496 23783 32548 23792
rect 32496 23749 32505 23783
rect 32505 23749 32539 23783
rect 32539 23749 32548 23783
rect 32496 23740 32548 23749
rect 34152 23783 34204 23792
rect 34152 23749 34161 23783
rect 34161 23749 34195 23783
rect 34195 23749 34204 23783
rect 34152 23740 34204 23749
rect 19616 23672 19668 23724
rect 19984 23672 20036 23724
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 29736 23647 29788 23656
rect 29736 23613 29745 23647
rect 29745 23613 29779 23647
rect 29779 23613 29788 23647
rect 29736 23604 29788 23613
rect 19340 23511 19392 23520
rect 19340 23477 19349 23511
rect 19349 23477 19383 23511
rect 19383 23477 19392 23511
rect 19340 23468 19392 23477
rect 20720 23468 20772 23520
rect 29184 23536 29236 23588
rect 32036 23468 32088 23520
rect 5174 23366 5226 23418
rect 5238 23366 5290 23418
rect 5302 23366 5354 23418
rect 5366 23366 5418 23418
rect 5430 23366 5482 23418
rect 13622 23366 13674 23418
rect 13686 23366 13738 23418
rect 13750 23366 13802 23418
rect 13814 23366 13866 23418
rect 13878 23366 13930 23418
rect 22070 23366 22122 23418
rect 22134 23366 22186 23418
rect 22198 23366 22250 23418
rect 22262 23366 22314 23418
rect 22326 23366 22378 23418
rect 30518 23366 30570 23418
rect 30582 23366 30634 23418
rect 30646 23366 30698 23418
rect 30710 23366 30762 23418
rect 30774 23366 30826 23418
rect 29736 23264 29788 23316
rect 30932 23196 30984 23248
rect 32680 23171 32732 23180
rect 32680 23137 32689 23171
rect 32689 23137 32723 23171
rect 32723 23137 32732 23171
rect 32680 23128 32732 23137
rect 19984 23103 20036 23112
rect 19984 23069 19993 23103
rect 19993 23069 20027 23103
rect 20027 23069 20036 23103
rect 19984 23060 20036 23069
rect 33140 23103 33192 23112
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 30840 22992 30892 23044
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 32496 22924 32548 22976
rect 9398 22822 9450 22874
rect 9462 22822 9514 22874
rect 9526 22822 9578 22874
rect 9590 22822 9642 22874
rect 9654 22822 9706 22874
rect 17846 22822 17898 22874
rect 17910 22822 17962 22874
rect 17974 22822 18026 22874
rect 18038 22822 18090 22874
rect 18102 22822 18154 22874
rect 26294 22822 26346 22874
rect 26358 22822 26410 22874
rect 26422 22822 26474 22874
rect 26486 22822 26538 22874
rect 26550 22822 26602 22874
rect 30840 22763 30892 22772
rect 30840 22729 30849 22763
rect 30849 22729 30883 22763
rect 30883 22729 30892 22763
rect 30840 22720 30892 22729
rect 32496 22695 32548 22704
rect 32496 22661 32505 22695
rect 32505 22661 32539 22695
rect 32539 22661 32548 22695
rect 32496 22652 32548 22661
rect 34152 22695 34204 22704
rect 34152 22661 34161 22695
rect 34161 22661 34195 22695
rect 34195 22661 34204 22695
rect 34152 22652 34204 22661
rect 30380 22584 30432 22636
rect 31116 22584 31168 22636
rect 32772 22516 32824 22568
rect 5174 22278 5226 22330
rect 5238 22278 5290 22330
rect 5302 22278 5354 22330
rect 5366 22278 5418 22330
rect 5430 22278 5482 22330
rect 13622 22278 13674 22330
rect 13686 22278 13738 22330
rect 13750 22278 13802 22330
rect 13814 22278 13866 22330
rect 13878 22278 13930 22330
rect 22070 22278 22122 22330
rect 22134 22278 22186 22330
rect 22198 22278 22250 22330
rect 22262 22278 22314 22330
rect 22326 22278 22378 22330
rect 30518 22278 30570 22330
rect 30582 22278 30634 22330
rect 30646 22278 30698 22330
rect 30710 22278 30762 22330
rect 30774 22278 30826 22330
rect 9398 21734 9450 21786
rect 9462 21734 9514 21786
rect 9526 21734 9578 21786
rect 9590 21734 9642 21786
rect 9654 21734 9706 21786
rect 17846 21734 17898 21786
rect 17910 21734 17962 21786
rect 17974 21734 18026 21786
rect 18038 21734 18090 21786
rect 18102 21734 18154 21786
rect 26294 21734 26346 21786
rect 26358 21734 26410 21786
rect 26422 21734 26474 21786
rect 26486 21734 26538 21786
rect 26550 21734 26602 21786
rect 17684 21539 17736 21548
rect 17684 21505 17693 21539
rect 17693 21505 17727 21539
rect 17727 21505 17736 21539
rect 17684 21496 17736 21505
rect 16948 21428 17000 21480
rect 23480 21428 23532 21480
rect 5174 21190 5226 21242
rect 5238 21190 5290 21242
rect 5302 21190 5354 21242
rect 5366 21190 5418 21242
rect 5430 21190 5482 21242
rect 13622 21190 13674 21242
rect 13686 21190 13738 21242
rect 13750 21190 13802 21242
rect 13814 21190 13866 21242
rect 13878 21190 13930 21242
rect 22070 21190 22122 21242
rect 22134 21190 22186 21242
rect 22198 21190 22250 21242
rect 22262 21190 22314 21242
rect 22326 21190 22378 21242
rect 30518 21190 30570 21242
rect 30582 21190 30634 21242
rect 30646 21190 30698 21242
rect 30710 21190 30762 21242
rect 30774 21190 30826 21242
rect 17224 20884 17276 20936
rect 17684 20884 17736 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 17592 20791 17644 20800
rect 17592 20757 17601 20791
rect 17601 20757 17635 20791
rect 17635 20757 17644 20791
rect 17592 20748 17644 20757
rect 9398 20646 9450 20698
rect 9462 20646 9514 20698
rect 9526 20646 9578 20698
rect 9590 20646 9642 20698
rect 9654 20646 9706 20698
rect 17846 20646 17898 20698
rect 17910 20646 17962 20698
rect 17974 20646 18026 20698
rect 18038 20646 18090 20698
rect 18102 20646 18154 20698
rect 26294 20646 26346 20698
rect 26358 20646 26410 20698
rect 26422 20646 26474 20698
rect 26486 20646 26538 20698
rect 26550 20646 26602 20698
rect 10324 20476 10376 20528
rect 16580 20408 16632 20460
rect 17040 20408 17092 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 32956 20476 33008 20528
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 20720 20408 20772 20460
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 29092 20272 29144 20324
rect 8484 20204 8536 20256
rect 8668 20204 8720 20256
rect 16856 20204 16908 20256
rect 24584 20204 24636 20256
rect 5174 20102 5226 20154
rect 5238 20102 5290 20154
rect 5302 20102 5354 20154
rect 5366 20102 5418 20154
rect 5430 20102 5482 20154
rect 13622 20102 13674 20154
rect 13686 20102 13738 20154
rect 13750 20102 13802 20154
rect 13814 20102 13866 20154
rect 13878 20102 13930 20154
rect 22070 20102 22122 20154
rect 22134 20102 22186 20154
rect 22198 20102 22250 20154
rect 22262 20102 22314 20154
rect 22326 20102 22378 20154
rect 30518 20102 30570 20154
rect 30582 20102 30634 20154
rect 30646 20102 30698 20154
rect 30710 20102 30762 20154
rect 30774 20102 30826 20154
rect 16304 20043 16356 20052
rect 16304 20009 16313 20043
rect 16313 20009 16347 20043
rect 16347 20009 16356 20043
rect 16304 20000 16356 20009
rect 17592 19932 17644 19984
rect 3516 19728 3568 19780
rect 17040 19907 17092 19916
rect 17040 19873 17049 19907
rect 17049 19873 17083 19907
rect 17083 19873 17092 19907
rect 17040 19864 17092 19873
rect 24584 19907 24636 19916
rect 24584 19873 24593 19907
rect 24593 19873 24627 19907
rect 24627 19873 24636 19907
rect 24584 19864 24636 19873
rect 9128 19796 9180 19848
rect 17408 19796 17460 19848
rect 29552 19907 29604 19916
rect 29552 19873 29561 19907
rect 29561 19873 29595 19907
rect 29595 19873 29604 19907
rect 29552 19864 29604 19873
rect 11612 19728 11664 19780
rect 16856 19728 16908 19780
rect 24308 19728 24360 19780
rect 31392 19771 31444 19780
rect 31392 19737 31401 19771
rect 31401 19737 31435 19771
rect 31435 19737 31444 19771
rect 31392 19728 31444 19737
rect 31760 19660 31812 19712
rect 9398 19558 9450 19610
rect 9462 19558 9514 19610
rect 9526 19558 9578 19610
rect 9590 19558 9642 19610
rect 9654 19558 9706 19610
rect 17846 19558 17898 19610
rect 17910 19558 17962 19610
rect 17974 19558 18026 19610
rect 18038 19558 18090 19610
rect 18102 19558 18154 19610
rect 26294 19558 26346 19610
rect 26358 19558 26410 19610
rect 26422 19558 26474 19610
rect 26486 19558 26538 19610
rect 26550 19558 26602 19610
rect 11612 19499 11664 19508
rect 11612 19465 11621 19499
rect 11621 19465 11655 19499
rect 11655 19465 11664 19499
rect 11612 19456 11664 19465
rect 8668 19431 8720 19440
rect 8668 19397 8677 19431
rect 8677 19397 8711 19431
rect 8711 19397 8720 19431
rect 8668 19388 8720 19397
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 10324 19363 10376 19372
rect 10324 19329 10333 19363
rect 10333 19329 10367 19363
rect 10367 19329 10376 19363
rect 10324 19320 10376 19329
rect 17132 19388 17184 19440
rect 20168 19456 20220 19508
rect 24308 19499 24360 19508
rect 24308 19465 24317 19499
rect 24317 19465 24351 19499
rect 24351 19465 24360 19499
rect 24308 19456 24360 19465
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17040 19252 17092 19304
rect 18236 19388 18288 19440
rect 18880 19388 18932 19440
rect 30380 19388 30432 19440
rect 17408 19320 17460 19372
rect 18696 19363 18748 19372
rect 17500 19184 17552 19236
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 23480 19320 23532 19372
rect 33048 19295 33100 19304
rect 33048 19261 33057 19295
rect 33057 19261 33091 19295
rect 33091 19261 33100 19295
rect 33048 19252 33100 19261
rect 33232 19252 33284 19304
rect 34152 19295 34204 19304
rect 34152 19261 34161 19295
rect 34161 19261 34195 19295
rect 34195 19261 34204 19295
rect 34152 19252 34204 19261
rect 6276 19116 6328 19168
rect 10232 19116 10284 19168
rect 5174 19014 5226 19066
rect 5238 19014 5290 19066
rect 5302 19014 5354 19066
rect 5366 19014 5418 19066
rect 5430 19014 5482 19066
rect 13622 19014 13674 19066
rect 13686 19014 13738 19066
rect 13750 19014 13802 19066
rect 13814 19014 13866 19066
rect 13878 19014 13930 19066
rect 22070 19014 22122 19066
rect 22134 19014 22186 19066
rect 22198 19014 22250 19066
rect 22262 19014 22314 19066
rect 22326 19014 22378 19066
rect 30518 19014 30570 19066
rect 30582 19014 30634 19066
rect 30646 19014 30698 19066
rect 30710 19014 30762 19066
rect 30774 19014 30826 19066
rect 9312 18912 9364 18964
rect 17316 18912 17368 18964
rect 17684 18912 17736 18964
rect 33232 18955 33284 18964
rect 33232 18921 33241 18955
rect 33241 18921 33275 18955
rect 33275 18921 33284 18955
rect 33232 18912 33284 18921
rect 34152 18912 34204 18964
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 5080 18708 5132 18760
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 10692 18819 10744 18828
rect 10692 18785 10701 18819
rect 10701 18785 10735 18819
rect 10735 18785 10744 18819
rect 10692 18776 10744 18785
rect 19156 18844 19208 18896
rect 19340 18776 19392 18828
rect 31668 18844 31720 18896
rect 9312 18708 9364 18760
rect 17224 18708 17276 18760
rect 27160 18751 27212 18760
rect 27160 18717 27169 18751
rect 27169 18717 27203 18751
rect 27203 18717 27212 18751
rect 27160 18708 27212 18717
rect 32036 18708 32088 18760
rect 32128 18708 32180 18760
rect 6644 18640 6696 18692
rect 8116 18683 8168 18692
rect 8116 18649 8125 18683
rect 8125 18649 8159 18683
rect 8159 18649 8168 18683
rect 8116 18640 8168 18649
rect 3424 18572 3476 18624
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 17408 18683 17460 18692
rect 17408 18649 17417 18683
rect 17417 18649 17451 18683
rect 17451 18649 17460 18683
rect 17408 18640 17460 18649
rect 27344 18683 27396 18692
rect 27344 18649 27353 18683
rect 27353 18649 27387 18683
rect 27387 18649 27396 18683
rect 27344 18640 27396 18649
rect 33324 18708 33376 18760
rect 33784 18708 33836 18760
rect 9036 18572 9088 18581
rect 10692 18572 10744 18624
rect 11060 18572 11112 18624
rect 16488 18615 16540 18624
rect 16488 18581 16497 18615
rect 16497 18581 16531 18615
rect 16531 18581 16540 18615
rect 16488 18572 16540 18581
rect 17776 18572 17828 18624
rect 32312 18572 32364 18624
rect 9398 18470 9450 18522
rect 9462 18470 9514 18522
rect 9526 18470 9578 18522
rect 9590 18470 9642 18522
rect 9654 18470 9706 18522
rect 17846 18470 17898 18522
rect 17910 18470 17962 18522
rect 17974 18470 18026 18522
rect 18038 18470 18090 18522
rect 18102 18470 18154 18522
rect 26294 18470 26346 18522
rect 26358 18470 26410 18522
rect 26422 18470 26474 18522
rect 26486 18470 26538 18522
rect 26550 18470 26602 18522
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 6736 18368 6788 18420
rect 16948 18368 17000 18420
rect 3424 18164 3476 18216
rect 17224 18300 17276 18352
rect 17592 18300 17644 18352
rect 32312 18343 32364 18352
rect 32312 18309 32321 18343
rect 32321 18309 32355 18343
rect 32355 18309 32364 18343
rect 32312 18300 32364 18309
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 9128 18275 9180 18284
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 17500 18232 17552 18284
rect 27160 18232 27212 18284
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 33876 18207 33928 18216
rect 6552 18028 6604 18080
rect 8484 18028 8536 18080
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 9036 18096 9088 18148
rect 33876 18173 33885 18207
rect 33885 18173 33919 18207
rect 33919 18173 33928 18207
rect 33876 18164 33928 18173
rect 17132 18071 17184 18080
rect 17132 18037 17141 18071
rect 17141 18037 17175 18071
rect 17175 18037 17184 18071
rect 17132 18028 17184 18037
rect 27160 18028 27212 18080
rect 29552 18071 29604 18080
rect 29552 18037 29561 18071
rect 29561 18037 29595 18071
rect 29595 18037 29604 18071
rect 29552 18028 29604 18037
rect 5174 17926 5226 17978
rect 5238 17926 5290 17978
rect 5302 17926 5354 17978
rect 5366 17926 5418 17978
rect 5430 17926 5482 17978
rect 13622 17926 13674 17978
rect 13686 17926 13738 17978
rect 13750 17926 13802 17978
rect 13814 17926 13866 17978
rect 13878 17926 13930 17978
rect 22070 17926 22122 17978
rect 22134 17926 22186 17978
rect 22198 17926 22250 17978
rect 22262 17926 22314 17978
rect 22326 17926 22378 17978
rect 30518 17926 30570 17978
rect 30582 17926 30634 17978
rect 30646 17926 30698 17978
rect 30710 17926 30762 17978
rect 30774 17926 30826 17978
rect 27344 17824 27396 17876
rect 6920 17756 6972 17808
rect 5080 17688 5132 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 8668 17688 8720 17740
rect 27804 17688 27856 17740
rect 29552 17731 29604 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 27160 17663 27212 17672
rect 27160 17629 27169 17663
rect 27169 17629 27203 17663
rect 27203 17629 27212 17663
rect 27160 17620 27212 17629
rect 28264 17620 28316 17672
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 33048 17688 33100 17740
rect 5356 17595 5408 17604
rect 5356 17561 5365 17595
rect 5365 17561 5399 17595
rect 5399 17561 5408 17595
rect 5356 17552 5408 17561
rect 8484 17552 8536 17604
rect 1584 17484 1636 17536
rect 7380 17484 7432 17536
rect 7840 17484 7892 17536
rect 25228 17484 25280 17536
rect 27712 17484 27764 17536
rect 9398 17382 9450 17434
rect 9462 17382 9514 17434
rect 9526 17382 9578 17434
rect 9590 17382 9642 17434
rect 9654 17382 9706 17434
rect 17846 17382 17898 17434
rect 17910 17382 17962 17434
rect 17974 17382 18026 17434
rect 18038 17382 18090 17434
rect 18102 17382 18154 17434
rect 26294 17382 26346 17434
rect 26358 17382 26410 17434
rect 26422 17382 26474 17434
rect 26486 17382 26538 17434
rect 26550 17382 26602 17434
rect 2044 17280 2096 17332
rect 5356 17323 5408 17332
rect 3056 17212 3108 17264
rect 5356 17289 5365 17323
rect 5365 17289 5399 17323
rect 5399 17289 5408 17323
rect 5356 17280 5408 17289
rect 27712 17255 27764 17264
rect 2780 17187 2832 17196
rect 2780 17153 2789 17187
rect 2789 17153 2823 17187
rect 2823 17153 2832 17187
rect 2780 17144 2832 17153
rect 27712 17221 27721 17255
rect 27721 17221 27755 17255
rect 27755 17221 27764 17255
rect 27712 17212 27764 17221
rect 3332 17119 3384 17128
rect 3332 17085 3341 17119
rect 3341 17085 3375 17119
rect 3375 17085 3384 17119
rect 3332 17076 3384 17085
rect 27528 17119 27580 17128
rect 27528 17085 27537 17119
rect 27537 17085 27571 17119
rect 27571 17085 27580 17119
rect 27528 17076 27580 17085
rect 32312 17076 32364 17128
rect 1400 16940 1452 16992
rect 32312 16940 32364 16992
rect 5174 16838 5226 16890
rect 5238 16838 5290 16890
rect 5302 16838 5354 16890
rect 5366 16838 5418 16890
rect 5430 16838 5482 16890
rect 13622 16838 13674 16890
rect 13686 16838 13738 16890
rect 13750 16838 13802 16890
rect 13814 16838 13866 16890
rect 13878 16838 13930 16890
rect 22070 16838 22122 16890
rect 22134 16838 22186 16890
rect 22198 16838 22250 16890
rect 22262 16838 22314 16890
rect 22326 16838 22378 16890
rect 30518 16838 30570 16890
rect 30582 16838 30634 16890
rect 30646 16838 30698 16890
rect 30710 16838 30762 16890
rect 30774 16838 30826 16890
rect 27528 16736 27580 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 32312 16643 32364 16652
rect 32312 16609 32321 16643
rect 32321 16609 32355 16643
rect 32355 16609 32364 16643
rect 32312 16600 32364 16609
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 32772 16464 32824 16516
rect 34152 16507 34204 16516
rect 34152 16473 34161 16507
rect 34161 16473 34195 16507
rect 34195 16473 34204 16507
rect 34152 16464 34204 16473
rect 9398 16294 9450 16346
rect 9462 16294 9514 16346
rect 9526 16294 9578 16346
rect 9590 16294 9642 16346
rect 9654 16294 9706 16346
rect 17846 16294 17898 16346
rect 17910 16294 17962 16346
rect 17974 16294 18026 16346
rect 18038 16294 18090 16346
rect 18102 16294 18154 16346
rect 26294 16294 26346 16346
rect 26358 16294 26410 16346
rect 26422 16294 26474 16346
rect 26486 16294 26538 16346
rect 26550 16294 26602 16346
rect 32772 16235 32824 16244
rect 32772 16201 32781 16235
rect 32781 16201 32815 16235
rect 32815 16201 32824 16235
rect 32772 16192 32824 16201
rect 17408 16167 17460 16176
rect 17408 16133 17417 16167
rect 17417 16133 17451 16167
rect 17451 16133 17460 16167
rect 17408 16124 17460 16133
rect 18236 16124 18288 16176
rect 33140 16124 33192 16176
rect 20812 15920 20864 15972
rect 32404 15988 32456 16040
rect 4252 15895 4304 15904
rect 4252 15861 4261 15895
rect 4261 15861 4295 15895
rect 4295 15861 4304 15895
rect 4252 15852 4304 15861
rect 8944 15852 8996 15904
rect 9128 15852 9180 15904
rect 16948 15852 17000 15904
rect 5174 15750 5226 15802
rect 5238 15750 5290 15802
rect 5302 15750 5354 15802
rect 5366 15750 5418 15802
rect 5430 15750 5482 15802
rect 13622 15750 13674 15802
rect 13686 15750 13738 15802
rect 13750 15750 13802 15802
rect 13814 15750 13866 15802
rect 13878 15750 13930 15802
rect 22070 15750 22122 15802
rect 22134 15750 22186 15802
rect 22198 15750 22250 15802
rect 22262 15750 22314 15802
rect 22326 15750 22378 15802
rect 30518 15750 30570 15802
rect 30582 15750 30634 15802
rect 30646 15750 30698 15802
rect 30710 15750 30762 15802
rect 30774 15750 30826 15802
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 4068 15580 4120 15632
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 9864 15555 9916 15564
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 17408 15444 17460 15496
rect 18972 15444 19024 15496
rect 20996 15444 21048 15496
rect 4436 15419 4488 15428
rect 4436 15385 4445 15419
rect 4445 15385 4479 15419
rect 4479 15385 4488 15419
rect 4436 15376 4488 15385
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 18972 15308 19024 15360
rect 9398 15206 9450 15258
rect 9462 15206 9514 15258
rect 9526 15206 9578 15258
rect 9590 15206 9642 15258
rect 9654 15206 9706 15258
rect 17846 15206 17898 15258
rect 17910 15206 17962 15258
rect 17974 15206 18026 15258
rect 18038 15206 18090 15258
rect 18102 15206 18154 15258
rect 26294 15206 26346 15258
rect 26358 15206 26410 15258
rect 26422 15206 26474 15258
rect 26486 15206 26538 15258
rect 26550 15206 26602 15258
rect 4436 15104 4488 15156
rect 10232 15104 10284 15156
rect 17500 15104 17552 15156
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 5632 14968 5684 15020
rect 18972 14968 19024 15020
rect 27160 14968 27212 15020
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 31024 14900 31076 14952
rect 31944 14900 31996 14952
rect 1584 14764 1636 14816
rect 25504 14764 25556 14816
rect 5174 14662 5226 14714
rect 5238 14662 5290 14714
rect 5302 14662 5354 14714
rect 5366 14662 5418 14714
rect 5430 14662 5482 14714
rect 13622 14662 13674 14714
rect 13686 14662 13738 14714
rect 13750 14662 13802 14714
rect 13814 14662 13866 14714
rect 13878 14662 13930 14714
rect 22070 14662 22122 14714
rect 22134 14662 22186 14714
rect 22198 14662 22250 14714
rect 22262 14662 22314 14714
rect 22326 14662 22378 14714
rect 30518 14662 30570 14714
rect 30582 14662 30634 14714
rect 30646 14662 30698 14714
rect 30710 14662 30762 14714
rect 30774 14662 30826 14714
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 25504 14467 25556 14476
rect 25504 14433 25513 14467
rect 25513 14433 25547 14467
rect 25547 14433 25556 14467
rect 25504 14424 25556 14433
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 25320 14399 25372 14408
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 31760 14288 31812 14340
rect 9398 14118 9450 14170
rect 9462 14118 9514 14170
rect 9526 14118 9578 14170
rect 9590 14118 9642 14170
rect 9654 14118 9706 14170
rect 17846 14118 17898 14170
rect 17910 14118 17962 14170
rect 17974 14118 18026 14170
rect 18038 14118 18090 14170
rect 18102 14118 18154 14170
rect 26294 14118 26346 14170
rect 26358 14118 26410 14170
rect 26422 14118 26474 14170
rect 26486 14118 26538 14170
rect 26550 14118 26602 14170
rect 1400 13880 1452 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 17684 13923 17736 13932
rect 17684 13889 17693 13923
rect 17693 13889 17727 13923
rect 17727 13889 17736 13923
rect 17684 13880 17736 13889
rect 25320 13923 25372 13932
rect 25320 13889 25329 13923
rect 25329 13889 25363 13923
rect 25363 13889 25372 13923
rect 25320 13880 25372 13889
rect 6184 13812 6236 13864
rect 6920 13812 6972 13864
rect 16856 13719 16908 13728
rect 16856 13685 16865 13719
rect 16865 13685 16899 13719
rect 16899 13685 16908 13719
rect 16856 13676 16908 13685
rect 17040 13676 17092 13728
rect 25964 13719 26016 13728
rect 25964 13685 25973 13719
rect 25973 13685 26007 13719
rect 26007 13685 26016 13719
rect 25964 13676 26016 13685
rect 32312 13676 32364 13728
rect 33968 13719 34020 13728
rect 33968 13685 33977 13719
rect 33977 13685 34011 13719
rect 34011 13685 34020 13719
rect 33968 13676 34020 13685
rect 5174 13574 5226 13626
rect 5238 13574 5290 13626
rect 5302 13574 5354 13626
rect 5366 13574 5418 13626
rect 5430 13574 5482 13626
rect 13622 13574 13674 13626
rect 13686 13574 13738 13626
rect 13750 13574 13802 13626
rect 13814 13574 13866 13626
rect 13878 13574 13930 13626
rect 22070 13574 22122 13626
rect 22134 13574 22186 13626
rect 22198 13574 22250 13626
rect 22262 13574 22314 13626
rect 22326 13574 22378 13626
rect 30518 13574 30570 13626
rect 30582 13574 30634 13626
rect 30646 13574 30698 13626
rect 30710 13574 30762 13626
rect 30774 13574 30826 13626
rect 6184 13404 6236 13456
rect 2780 13336 2832 13388
rect 16764 13404 16816 13456
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 25964 13336 26016 13388
rect 32772 13336 32824 13388
rect 33048 13379 33100 13388
rect 33048 13345 33057 13379
rect 33057 13345 33091 13379
rect 33091 13345 33100 13379
rect 33048 13336 33100 13345
rect 33968 13336 34020 13388
rect 8208 13268 8260 13320
rect 9956 13268 10008 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 6920 13243 6972 13252
rect 6920 13209 6929 13243
rect 6929 13209 6963 13243
rect 6963 13209 6972 13243
rect 25596 13243 25648 13252
rect 6920 13200 6972 13209
rect 25596 13209 25605 13243
rect 25605 13209 25639 13243
rect 25639 13209 25648 13243
rect 25596 13200 25648 13209
rect 33968 13243 34020 13252
rect 33968 13209 33977 13243
rect 33977 13209 34011 13243
rect 34011 13209 34020 13243
rect 33968 13200 34020 13209
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 9398 13030 9450 13082
rect 9462 13030 9514 13082
rect 9526 13030 9578 13082
rect 9590 13030 9642 13082
rect 9654 13030 9706 13082
rect 17846 13030 17898 13082
rect 17910 13030 17962 13082
rect 17974 13030 18026 13082
rect 18038 13030 18090 13082
rect 18102 13030 18154 13082
rect 26294 13030 26346 13082
rect 26358 13030 26410 13082
rect 26422 13030 26474 13082
rect 26486 13030 26538 13082
rect 26550 13030 26602 13082
rect 5632 12928 5684 12980
rect 14372 12928 14424 12980
rect 25596 12928 25648 12980
rect 34152 12903 34204 12912
rect 34152 12869 34161 12903
rect 34161 12869 34195 12903
rect 34195 12869 34204 12903
rect 34152 12860 34204 12869
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 25320 12835 25372 12844
rect 8208 12792 8260 12801
rect 25320 12801 25329 12835
rect 25329 12801 25363 12835
rect 25363 12801 25372 12835
rect 25320 12792 25372 12801
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 4160 12724 4212 12776
rect 32496 12767 32548 12776
rect 32496 12733 32505 12767
rect 32505 12733 32539 12767
rect 32539 12733 32548 12767
rect 32496 12724 32548 12733
rect 14372 12588 14424 12640
rect 16304 12588 16356 12640
rect 5174 12486 5226 12538
rect 5238 12486 5290 12538
rect 5302 12486 5354 12538
rect 5366 12486 5418 12538
rect 5430 12486 5482 12538
rect 13622 12486 13674 12538
rect 13686 12486 13738 12538
rect 13750 12486 13802 12538
rect 13814 12486 13866 12538
rect 13878 12486 13930 12538
rect 22070 12486 22122 12538
rect 22134 12486 22186 12538
rect 22198 12486 22250 12538
rect 22262 12486 22314 12538
rect 22326 12486 22378 12538
rect 30518 12486 30570 12538
rect 30582 12486 30634 12538
rect 30646 12486 30698 12538
rect 30710 12486 30762 12538
rect 30774 12486 30826 12538
rect 32496 12384 32548 12436
rect 33968 12384 34020 12436
rect 32496 12223 32548 12232
rect 32496 12189 32505 12223
rect 32505 12189 32539 12223
rect 32539 12189 32548 12223
rect 32496 12180 32548 12189
rect 33784 12223 33836 12232
rect 33784 12189 33793 12223
rect 33793 12189 33827 12223
rect 33827 12189 33836 12223
rect 33784 12180 33836 12189
rect 9398 11942 9450 11994
rect 9462 11942 9514 11994
rect 9526 11942 9578 11994
rect 9590 11942 9642 11994
rect 9654 11942 9706 11994
rect 17846 11942 17898 11994
rect 17910 11942 17962 11994
rect 17974 11942 18026 11994
rect 18038 11942 18090 11994
rect 18102 11942 18154 11994
rect 26294 11942 26346 11994
rect 26358 11942 26410 11994
rect 26422 11942 26474 11994
rect 26486 11942 26538 11994
rect 26550 11942 26602 11994
rect 17776 11704 17828 11756
rect 20812 11704 20864 11756
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 16856 11500 16908 11552
rect 17040 11500 17092 11552
rect 20904 11500 20956 11552
rect 5174 11398 5226 11450
rect 5238 11398 5290 11450
rect 5302 11398 5354 11450
rect 5366 11398 5418 11450
rect 5430 11398 5482 11450
rect 13622 11398 13674 11450
rect 13686 11398 13738 11450
rect 13750 11398 13802 11450
rect 13814 11398 13866 11450
rect 13878 11398 13930 11450
rect 22070 11398 22122 11450
rect 22134 11398 22186 11450
rect 22198 11398 22250 11450
rect 22262 11398 22314 11450
rect 22326 11398 22378 11450
rect 30518 11398 30570 11450
rect 30582 11398 30634 11450
rect 30646 11398 30698 11450
rect 30710 11398 30762 11450
rect 30774 11398 30826 11450
rect 664 11160 716 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 21732 11203 21784 11212
rect 21732 11169 21741 11203
rect 21741 11169 21775 11203
rect 21775 11169 21784 11203
rect 21732 11160 21784 11169
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 9128 11092 9180 11144
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 3332 11024 3384 11076
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 9398 10854 9450 10906
rect 9462 10854 9514 10906
rect 9526 10854 9578 10906
rect 9590 10854 9642 10906
rect 9654 10854 9706 10906
rect 17846 10854 17898 10906
rect 17910 10854 17962 10906
rect 17974 10854 18026 10906
rect 18038 10854 18090 10906
rect 18102 10854 18154 10906
rect 26294 10854 26346 10906
rect 26358 10854 26410 10906
rect 26422 10854 26474 10906
rect 26486 10854 26538 10906
rect 26550 10854 26602 10906
rect 7104 10752 7156 10804
rect 14464 10795 14516 10804
rect 14464 10761 14473 10795
rect 14473 10761 14507 10795
rect 14507 10761 14516 10795
rect 14464 10752 14516 10761
rect 2872 10684 2924 10736
rect 2320 10616 2372 10668
rect 17684 10684 17736 10736
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 27068 10616 27120 10668
rect 2780 10548 2832 10600
rect 7288 10548 7340 10600
rect 9772 10548 9824 10600
rect 27804 10591 27856 10600
rect 8944 10480 8996 10532
rect 27804 10557 27813 10591
rect 27813 10557 27847 10591
rect 27847 10557 27856 10591
rect 27804 10548 27856 10557
rect 31668 10548 31720 10600
rect 5174 10310 5226 10362
rect 5238 10310 5290 10362
rect 5302 10310 5354 10362
rect 5366 10310 5418 10362
rect 5430 10310 5482 10362
rect 13622 10310 13674 10362
rect 13686 10310 13738 10362
rect 13750 10310 13802 10362
rect 13814 10310 13866 10362
rect 13878 10310 13930 10362
rect 22070 10310 22122 10362
rect 22134 10310 22186 10362
rect 22198 10310 22250 10362
rect 22262 10310 22314 10362
rect 22326 10310 22378 10362
rect 30518 10310 30570 10362
rect 30582 10310 30634 10362
rect 30646 10310 30698 10362
rect 30710 10310 30762 10362
rect 30774 10310 30826 10362
rect 9772 10251 9824 10260
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 27804 10208 27856 10260
rect 1952 10072 2004 10124
rect 10416 10072 10468 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 2964 10004 3016 10056
rect 11888 10004 11940 10056
rect 16488 10004 16540 10056
rect 28264 10004 28316 10056
rect 12164 9936 12216 9988
rect 1584 9868 1636 9920
rect 2964 9911 3016 9920
rect 2964 9877 2973 9911
rect 2973 9877 3007 9911
rect 3007 9877 3016 9911
rect 2964 9868 3016 9877
rect 12072 9868 12124 9920
rect 16488 9868 16540 9920
rect 16672 9868 16724 9920
rect 19616 9911 19668 9920
rect 19616 9877 19625 9911
rect 19625 9877 19659 9911
rect 19659 9877 19668 9911
rect 19616 9868 19668 9877
rect 9398 9766 9450 9818
rect 9462 9766 9514 9818
rect 9526 9766 9578 9818
rect 9590 9766 9642 9818
rect 9654 9766 9706 9818
rect 17846 9766 17898 9818
rect 17910 9766 17962 9818
rect 17974 9766 18026 9818
rect 18038 9766 18090 9818
rect 18102 9766 18154 9818
rect 26294 9766 26346 9818
rect 26358 9766 26410 9818
rect 26422 9766 26474 9818
rect 26486 9766 26538 9818
rect 26550 9766 26602 9818
rect 2964 9596 3016 9648
rect 12072 9639 12124 9648
rect 12072 9605 12081 9639
rect 12081 9605 12115 9639
rect 12115 9605 12124 9639
rect 12072 9596 12124 9605
rect 12164 9596 12216 9648
rect 16488 9596 16540 9648
rect 19616 9639 19668 9648
rect 19616 9605 19625 9639
rect 19625 9605 19659 9639
rect 19659 9605 19668 9639
rect 19616 9596 19668 9605
rect 2412 9528 2464 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 2780 9460 2832 9512
rect 13452 9503 13504 9512
rect 13452 9469 13461 9503
rect 13461 9469 13495 9503
rect 13495 9469 13504 9503
rect 13452 9460 13504 9469
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 19984 9503 20036 9512
rect 19984 9469 19993 9503
rect 19993 9469 20027 9503
rect 20027 9469 20036 9503
rect 19984 9460 20036 9469
rect 1400 9324 1452 9376
rect 5174 9222 5226 9274
rect 5238 9222 5290 9274
rect 5302 9222 5354 9274
rect 5366 9222 5418 9274
rect 5430 9222 5482 9274
rect 13622 9222 13674 9274
rect 13686 9222 13738 9274
rect 13750 9222 13802 9274
rect 13814 9222 13866 9274
rect 13878 9222 13930 9274
rect 22070 9222 22122 9274
rect 22134 9222 22186 9274
rect 22198 9222 22250 9274
rect 22262 9222 22314 9274
rect 22326 9222 22378 9274
rect 30518 9222 30570 9274
rect 30582 9222 30634 9274
rect 30646 9222 30698 9274
rect 30710 9222 30762 9274
rect 30774 9222 30826 9274
rect 19432 9120 19484 9172
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 20812 8984 20864 9036
rect 23940 8916 23992 8968
rect 30932 8959 30984 8968
rect 30932 8925 30941 8959
rect 30941 8925 30975 8959
rect 30975 8925 30984 8959
rect 30932 8916 30984 8925
rect 30840 8848 30892 8900
rect 32772 8891 32824 8900
rect 32772 8857 32781 8891
rect 32781 8857 32815 8891
rect 32815 8857 32824 8891
rect 32772 8848 32824 8857
rect 24124 8780 24176 8832
rect 9398 8678 9450 8730
rect 9462 8678 9514 8730
rect 9526 8678 9578 8730
rect 9590 8678 9642 8730
rect 9654 8678 9706 8730
rect 17846 8678 17898 8730
rect 17910 8678 17962 8730
rect 17974 8678 18026 8730
rect 18038 8678 18090 8730
rect 18102 8678 18154 8730
rect 26294 8678 26346 8730
rect 26358 8678 26410 8730
rect 26422 8678 26474 8730
rect 26486 8678 26538 8730
rect 26550 8678 26602 8730
rect 30840 8619 30892 8628
rect 30840 8585 30849 8619
rect 30849 8585 30883 8619
rect 30883 8585 30892 8619
rect 30840 8576 30892 8585
rect 24124 8551 24176 8560
rect 24124 8517 24133 8551
rect 24133 8517 24167 8551
rect 24167 8517 24176 8551
rect 24124 8508 24176 8517
rect 12164 8440 12216 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 28264 8440 28316 8492
rect 31024 8508 31076 8560
rect 30932 8440 30984 8492
rect 12900 8372 12952 8424
rect 24492 8415 24544 8424
rect 24492 8381 24501 8415
rect 24501 8381 24535 8415
rect 24535 8381 24544 8415
rect 24492 8372 24544 8381
rect 13084 8304 13136 8356
rect 3148 8236 3200 8288
rect 9864 8236 9916 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 29736 8279 29788 8288
rect 29736 8245 29745 8279
rect 29745 8245 29779 8279
rect 29779 8245 29788 8279
rect 29736 8236 29788 8245
rect 5174 8134 5226 8186
rect 5238 8134 5290 8186
rect 5302 8134 5354 8186
rect 5366 8134 5418 8186
rect 5430 8134 5482 8186
rect 13622 8134 13674 8186
rect 13686 8134 13738 8186
rect 13750 8134 13802 8186
rect 13814 8134 13866 8186
rect 13878 8134 13930 8186
rect 22070 8134 22122 8186
rect 22134 8134 22186 8186
rect 22198 8134 22250 8186
rect 22262 8134 22314 8186
rect 22326 8134 22378 8186
rect 30518 8134 30570 8186
rect 30582 8134 30634 8186
rect 30646 8134 30698 8186
rect 30710 8134 30762 8186
rect 30774 8134 30826 8186
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 13084 7939 13136 7948
rect 13084 7905 13093 7939
rect 13093 7905 13127 7939
rect 13127 7905 13136 7939
rect 13084 7896 13136 7905
rect 29736 7896 29788 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 10048 7760 10100 7812
rect 29184 7760 29236 7812
rect 33048 7760 33100 7812
rect 9398 7590 9450 7642
rect 9462 7590 9514 7642
rect 9526 7590 9578 7642
rect 9590 7590 9642 7642
rect 9654 7590 9706 7642
rect 17846 7590 17898 7642
rect 17910 7590 17962 7642
rect 17974 7590 18026 7642
rect 18038 7590 18090 7642
rect 18102 7590 18154 7642
rect 26294 7590 26346 7642
rect 26358 7590 26410 7642
rect 26422 7590 26474 7642
rect 26486 7590 26538 7642
rect 26550 7590 26602 7642
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 6552 7352 6604 7404
rect 20996 7352 21048 7404
rect 2964 7284 3016 7336
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 7104 7148 7156 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 32680 7191 32732 7200
rect 32680 7157 32689 7191
rect 32689 7157 32723 7191
rect 32723 7157 32732 7191
rect 32680 7148 32732 7157
rect 5174 7046 5226 7098
rect 5238 7046 5290 7098
rect 5302 7046 5354 7098
rect 5366 7046 5418 7098
rect 5430 7046 5482 7098
rect 13622 7046 13674 7098
rect 13686 7046 13738 7098
rect 13750 7046 13802 7098
rect 13814 7046 13866 7098
rect 13878 7046 13930 7098
rect 22070 7046 22122 7098
rect 22134 7046 22186 7098
rect 22198 7046 22250 7098
rect 22262 7046 22314 7098
rect 22326 7046 22378 7098
rect 30518 7046 30570 7098
rect 30582 7046 30634 7098
rect 30646 7046 30698 7098
rect 30710 7046 30762 7098
rect 30774 7046 30826 7098
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 7288 6808 7340 6860
rect 20076 6851 20128 6860
rect 20076 6817 20085 6851
rect 20085 6817 20119 6851
rect 20119 6817 20128 6851
rect 20076 6808 20128 6817
rect 20812 6808 20864 6860
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10140 6740 10192 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 19708 6740 19760 6792
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 7104 6672 7156 6724
rect 20628 6672 20680 6724
rect 32680 6808 32732 6860
rect 34152 6851 34204 6860
rect 34152 6817 34161 6851
rect 34161 6817 34195 6851
rect 34195 6817 34204 6851
rect 34152 6808 34204 6817
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 30932 6740 30984 6792
rect 31208 6783 31260 6792
rect 31208 6749 31217 6783
rect 31217 6749 31251 6783
rect 31251 6749 31260 6783
rect 31208 6740 31260 6749
rect 32588 6672 32640 6724
rect 9772 6604 9824 6656
rect 12992 6604 13044 6656
rect 15752 6604 15804 6656
rect 30932 6604 30984 6656
rect 9398 6502 9450 6554
rect 9462 6502 9514 6554
rect 9526 6502 9578 6554
rect 9590 6502 9642 6554
rect 9654 6502 9706 6554
rect 17846 6502 17898 6554
rect 17910 6502 17962 6554
rect 17974 6502 18026 6554
rect 18038 6502 18090 6554
rect 18102 6502 18154 6554
rect 26294 6502 26346 6554
rect 26358 6502 26410 6554
rect 26422 6502 26474 6554
rect 26486 6502 26538 6554
rect 26550 6502 26602 6554
rect 18880 6400 18932 6452
rect 32588 6443 32640 6452
rect 32588 6409 32597 6443
rect 32597 6409 32631 6443
rect 32631 6409 32640 6443
rect 32588 6400 32640 6409
rect 12992 6375 13044 6384
rect 12992 6341 13001 6375
rect 13001 6341 13035 6375
rect 13035 6341 13044 6375
rect 12992 6332 13044 6341
rect 17132 6332 17184 6384
rect 32128 6332 32180 6384
rect 32404 6332 32456 6384
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 27252 6307 27304 6316
rect 27252 6273 27261 6307
rect 27261 6273 27295 6307
rect 27295 6273 27304 6307
rect 27252 6264 27304 6273
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 13268 6239 13320 6248
rect 5632 6128 5684 6180
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 26976 6196 27028 6248
rect 29092 6239 29144 6248
rect 29092 6205 29101 6239
rect 29101 6205 29135 6239
rect 29135 6205 29144 6239
rect 29092 6196 29144 6205
rect 10324 6060 10376 6112
rect 15936 6060 15988 6112
rect 5174 5958 5226 6010
rect 5238 5958 5290 6010
rect 5302 5958 5354 6010
rect 5366 5958 5418 6010
rect 5430 5958 5482 6010
rect 13622 5958 13674 6010
rect 13686 5958 13738 6010
rect 13750 5958 13802 6010
rect 13814 5958 13866 6010
rect 13878 5958 13930 6010
rect 22070 5958 22122 6010
rect 22134 5958 22186 6010
rect 22198 5958 22250 6010
rect 22262 5958 22314 6010
rect 22326 5958 22378 6010
rect 30518 5958 30570 6010
rect 30582 5958 30634 6010
rect 30646 5958 30698 6010
rect 30710 5958 30762 6010
rect 30774 5958 30826 6010
rect 26976 5899 27028 5908
rect 26976 5865 26985 5899
rect 26985 5865 27019 5899
rect 27019 5865 27028 5899
rect 26976 5856 27028 5865
rect 7104 5720 7156 5772
rect 10140 5763 10192 5772
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 31208 5788 31260 5840
rect 30932 5720 30984 5772
rect 32220 5763 32272 5772
rect 32220 5729 32229 5763
rect 32229 5729 32263 5763
rect 32263 5729 32272 5763
rect 32220 5720 32272 5729
rect 9036 5652 9088 5704
rect 19708 5652 19760 5704
rect 27620 5695 27672 5704
rect 27620 5661 27629 5695
rect 27629 5661 27663 5695
rect 27663 5661 27672 5695
rect 27620 5652 27672 5661
rect 7932 5584 7984 5636
rect 8392 5627 8444 5636
rect 8392 5593 8401 5627
rect 8401 5593 8435 5627
rect 8435 5593 8444 5627
rect 8392 5584 8444 5593
rect 13544 5584 13596 5636
rect 9398 5414 9450 5466
rect 9462 5414 9514 5466
rect 9526 5414 9578 5466
rect 9590 5414 9642 5466
rect 9654 5414 9706 5466
rect 17846 5414 17898 5466
rect 17910 5414 17962 5466
rect 17974 5414 18026 5466
rect 18038 5414 18090 5466
rect 18102 5414 18154 5466
rect 26294 5414 26346 5466
rect 26358 5414 26410 5466
rect 26422 5414 26474 5466
rect 26486 5414 26538 5466
rect 26550 5414 26602 5466
rect 8116 5312 8168 5364
rect 3424 5244 3476 5296
rect 10600 5312 10652 5364
rect 27620 5312 27672 5364
rect 9772 5244 9824 5296
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 17132 5176 17184 5228
rect 30380 5176 30432 5228
rect 10692 5108 10744 5160
rect 8208 5040 8260 5092
rect 27344 5108 27396 5160
rect 32312 5108 32364 5160
rect 29092 5040 29144 5092
rect 32404 5040 32456 5092
rect 7104 4972 7156 5024
rect 11152 4972 11204 5024
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 30380 5015 30432 5024
rect 30380 4981 30389 5015
rect 30389 4981 30423 5015
rect 30423 4981 30432 5015
rect 30380 4972 30432 4981
rect 5174 4870 5226 4922
rect 5238 4870 5290 4922
rect 5302 4870 5354 4922
rect 5366 4870 5418 4922
rect 5430 4870 5482 4922
rect 13622 4870 13674 4922
rect 13686 4870 13738 4922
rect 13750 4870 13802 4922
rect 13814 4870 13866 4922
rect 13878 4870 13930 4922
rect 22070 4870 22122 4922
rect 22134 4870 22186 4922
rect 22198 4870 22250 4922
rect 22262 4870 22314 4922
rect 22326 4870 22378 4922
rect 30518 4870 30570 4922
rect 30582 4870 30634 4922
rect 30646 4870 30698 4922
rect 30710 4870 30762 4922
rect 30774 4870 30826 4922
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 3424 4700 3476 4752
rect 13268 4768 13320 4820
rect 27344 4811 27396 4820
rect 27344 4777 27353 4811
rect 27353 4777 27387 4811
rect 27387 4777 27396 4811
rect 27344 4768 27396 4777
rect 6644 4632 6696 4684
rect 11612 4700 11664 4752
rect 30380 4700 30432 4752
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 7656 4564 7708 4616
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 30932 4632 30984 4641
rect 25320 4564 25372 4616
rect 30288 4607 30340 4616
rect 30288 4573 30297 4607
rect 30297 4573 30331 4607
rect 30331 4573 30340 4607
rect 30288 4564 30340 4573
rect 5540 4496 5592 4548
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 9398 4326 9450 4378
rect 9462 4326 9514 4378
rect 9526 4326 9578 4378
rect 9590 4326 9642 4378
rect 9654 4326 9706 4378
rect 17846 4326 17898 4378
rect 17910 4326 17962 4378
rect 17974 4326 18026 4378
rect 18038 4326 18090 4378
rect 18102 4326 18154 4378
rect 26294 4326 26346 4378
rect 26358 4326 26410 4378
rect 26422 4326 26474 4378
rect 26486 4326 26538 4378
rect 26550 4326 26602 4378
rect 7288 4199 7340 4208
rect 7288 4165 7297 4199
rect 7297 4165 7331 4199
rect 7331 4165 7340 4199
rect 7288 4156 7340 4165
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 30288 4131 30340 4140
rect 3424 4020 3476 4072
rect 3884 3952 3936 4004
rect 7656 4020 7708 4072
rect 30288 4097 30297 4131
rect 30297 4097 30331 4131
rect 30331 4097 30340 4131
rect 30288 4088 30340 4097
rect 32128 4088 32180 4140
rect 7840 3884 7892 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 32496 3884 32548 3936
rect 32864 3927 32916 3936
rect 32864 3893 32873 3927
rect 32873 3893 32907 3927
rect 32907 3893 32916 3927
rect 32864 3884 32916 3893
rect 5174 3782 5226 3834
rect 5238 3782 5290 3834
rect 5302 3782 5354 3834
rect 5366 3782 5418 3834
rect 5430 3782 5482 3834
rect 13622 3782 13674 3834
rect 13686 3782 13738 3834
rect 13750 3782 13802 3834
rect 13814 3782 13866 3834
rect 13878 3782 13930 3834
rect 22070 3782 22122 3834
rect 22134 3782 22186 3834
rect 22198 3782 22250 3834
rect 22262 3782 22314 3834
rect 22326 3782 22378 3834
rect 30518 3782 30570 3834
rect 30582 3782 30634 3834
rect 30646 3782 30698 3834
rect 30710 3782 30762 3834
rect 30774 3782 30826 3834
rect 5080 3544 5132 3596
rect 10232 3680 10284 3732
rect 10508 3612 10560 3664
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 9956 3544 10008 3553
rect 10324 3587 10376 3596
rect 10324 3553 10333 3587
rect 10333 3553 10367 3587
rect 10367 3553 10376 3587
rect 10324 3544 10376 3553
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 32864 3612 32916 3664
rect 32496 3587 32548 3596
rect 32496 3553 32505 3587
rect 32505 3553 32539 3587
rect 32539 3553 32548 3587
rect 32496 3544 32548 3553
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 17592 3476 17644 3528
rect 15752 3451 15804 3460
rect 15752 3417 15761 3451
rect 15761 3417 15795 3451
rect 15795 3417 15804 3451
rect 15752 3408 15804 3417
rect 34796 3408 34848 3460
rect 3240 3340 3292 3392
rect 6184 3340 6236 3392
rect 9398 3238 9450 3290
rect 9462 3238 9514 3290
rect 9526 3238 9578 3290
rect 9590 3238 9642 3290
rect 9654 3238 9706 3290
rect 17846 3238 17898 3290
rect 17910 3238 17962 3290
rect 17974 3238 18026 3290
rect 18038 3238 18090 3290
rect 18102 3238 18154 3290
rect 26294 3238 26346 3290
rect 26358 3238 26410 3290
rect 26422 3238 26474 3290
rect 26486 3238 26538 3290
rect 26550 3238 26602 3290
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 2596 2864 2648 2916
rect 35440 2932 35492 2984
rect 3424 2864 3476 2916
rect 8944 2864 8996 2916
rect 4528 2796 4580 2848
rect 5540 2796 5592 2848
rect 6460 2796 6512 2848
rect 8208 2796 8260 2848
rect 5174 2694 5226 2746
rect 5238 2694 5290 2746
rect 5302 2694 5354 2746
rect 5366 2694 5418 2746
rect 5430 2694 5482 2746
rect 13622 2694 13674 2746
rect 13686 2694 13738 2746
rect 13750 2694 13802 2746
rect 13814 2694 13866 2746
rect 13878 2694 13930 2746
rect 22070 2694 22122 2746
rect 22134 2694 22186 2746
rect 22198 2694 22250 2746
rect 22262 2694 22314 2746
rect 22326 2694 22378 2746
rect 30518 2694 30570 2746
rect 30582 2694 30634 2746
rect 30646 2694 30698 2746
rect 30710 2694 30762 2746
rect 30774 2694 30826 2746
rect 2964 2592 3016 2644
rect 15752 2635 15804 2644
rect 15752 2601 15761 2635
rect 15761 2601 15795 2635
rect 15795 2601 15804 2635
rect 15752 2592 15804 2601
rect 13452 2524 13504 2576
rect 31760 2592 31812 2644
rect 3056 2388 3108 2440
rect 16948 2388 17000 2440
rect 3424 2252 3476 2304
rect 5632 2252 5684 2304
rect 9398 2150 9450 2202
rect 9462 2150 9514 2202
rect 9526 2150 9578 2202
rect 9590 2150 9642 2202
rect 9654 2150 9706 2202
rect 17846 2150 17898 2202
rect 17910 2150 17962 2202
rect 17974 2150 18026 2202
rect 18038 2150 18090 2202
rect 18102 2150 18154 2202
rect 26294 2150 26346 2202
rect 26358 2150 26410 2202
rect 26422 2150 26474 2202
rect 26486 2150 26538 2202
rect 26550 2150 26602 2202
<< metal2 >>
rect -10 41200 102 42000
rect 634 41200 746 42000
rect 1278 41200 1390 42000
rect 1922 41200 2034 42000
rect 2566 41200 2678 42000
rect 3210 41200 3322 42000
rect 3606 41576 3662 41585
rect 3606 41511 3662 41520
rect 20 38548 72 38554
rect 20 38490 72 38496
rect 32 31278 60 38490
rect 676 37262 704 41200
rect 1320 38554 1348 41200
rect 1308 38548 1360 38554
rect 1308 38490 1360 38496
rect 3330 37496 3386 37505
rect 3330 37431 3386 37440
rect 664 37256 716 37262
rect 664 37198 716 37204
rect 1858 36136 1914 36145
rect 1858 36071 1860 36080
rect 1912 36071 1914 36080
rect 1860 36042 1912 36048
rect 1952 36032 2004 36038
rect 1952 35974 2004 35980
rect 20 31272 72 31278
rect 20 31214 72 31220
rect 1964 23730 1992 35974
rect 3344 35894 3372 37431
rect 3344 35866 3556 35894
rect 3330 35456 3386 35465
rect 3330 35391 3386 35400
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2792 30258 2820 30670
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 3148 30184 3200 30190
rect 3148 30126 3200 30132
rect 3160 29850 3188 30126
rect 3148 29844 3200 29850
rect 3148 29786 3200 29792
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2976 29306 3004 29582
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1596 16658 1624 17478
rect 2056 17338 2084 17614
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 2056 16574 2084 17274
rect 2792 17202 2820 17614
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 1964 16546 2084 16574
rect 1964 15026 1992 16546
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14482 1624 14758
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1400 14408 1452 14414
rect 1872 14385 1900 14418
rect 1400 14350 1452 14356
rect 1858 14376 1914 14385
rect 1412 13938 1440 14350
rect 1858 14311 1914 14320
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 664 11212 716 11218
rect 664 11154 716 11160
rect 676 800 704 11154
rect 1964 10130 1992 14962
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2792 13394 2820 13631
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2976 11150 3004 29242
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2332 10674 2360 11086
rect 2872 11008 2924 11014
rect 2778 10976 2834 10985
rect 2872 10950 2924 10956
rect 2778 10911 2834 10920
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2792 10606 2820 10911
rect 2884 10742 2912 10950
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2976 10062 3004 11086
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9042 1440 9318
rect 1596 9042 1624 9862
rect 2424 9586 2452 9998
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9654 3004 9862
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 8945 1900 8978
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7410 2452 7822
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2792 4865 2820 9454
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2976 6866 3004 7278
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3068 6798 3096 17206
rect 3344 17134 3372 35391
rect 3422 34096 3478 34105
rect 3422 34031 3478 34040
rect 3436 33930 3464 34031
rect 3424 33924 3476 33930
rect 3424 33866 3476 33872
rect 3422 32056 3478 32065
rect 3422 31991 3478 32000
rect 3436 31822 3464 31991
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3422 31376 3478 31385
rect 3422 31311 3478 31320
rect 3436 29578 3464 31311
rect 3424 29572 3476 29578
rect 3424 29514 3476 29520
rect 3422 25256 3478 25265
rect 3422 25191 3478 25200
rect 3436 24954 3464 25191
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3528 19786 3556 35866
rect 3620 25974 3648 41511
rect 4498 41200 4610 42000
rect 5142 41200 5254 42000
rect 5786 41200 5898 42000
rect 6012 41262 6316 41290
rect 5828 41154 5856 41200
rect 6012 41154 6040 41262
rect 5828 41126 6040 41154
rect 4066 40896 4122 40905
rect 4066 40831 4122 40840
rect 4080 38486 4108 40831
rect 5174 39740 5482 39749
rect 5174 39738 5180 39740
rect 5236 39738 5260 39740
rect 5316 39738 5340 39740
rect 5396 39738 5420 39740
rect 5476 39738 5482 39740
rect 5236 39686 5238 39738
rect 5418 39686 5420 39738
rect 5174 39684 5180 39686
rect 5236 39684 5260 39686
rect 5316 39684 5340 39686
rect 5396 39684 5420 39686
rect 5476 39684 5482 39686
rect 5174 39675 5482 39684
rect 4896 38752 4948 38758
rect 4896 38694 4948 38700
rect 4068 38480 4120 38486
rect 4068 38422 4120 38428
rect 4908 38418 4936 38694
rect 5174 38652 5482 38661
rect 5174 38650 5180 38652
rect 5236 38650 5260 38652
rect 5316 38650 5340 38652
rect 5396 38650 5420 38652
rect 5476 38650 5482 38652
rect 5236 38598 5238 38650
rect 5418 38598 5420 38650
rect 5174 38596 5180 38598
rect 5236 38596 5260 38598
rect 5316 38596 5340 38598
rect 5396 38596 5420 38598
rect 5476 38596 5482 38598
rect 5174 38587 5482 38596
rect 6288 38570 6316 41262
rect 6430 41200 6542 42000
rect 7074 41200 7186 42000
rect 7300 41262 7604 41290
rect 6288 38542 6868 38570
rect 4896 38412 4948 38418
rect 4896 38354 4948 38360
rect 6736 38344 6788 38350
rect 6736 38286 6788 38292
rect 5540 38276 5592 38282
rect 5540 38218 5592 38224
rect 5552 38010 5580 38218
rect 5540 38004 5592 38010
rect 5540 37946 5592 37952
rect 6748 37874 6776 38286
rect 6736 37868 6788 37874
rect 6736 37810 6788 37816
rect 5174 37564 5482 37573
rect 5174 37562 5180 37564
rect 5236 37562 5260 37564
rect 5316 37562 5340 37564
rect 5396 37562 5420 37564
rect 5476 37562 5482 37564
rect 5236 37510 5238 37562
rect 5418 37510 5420 37562
rect 5174 37508 5180 37510
rect 5236 37508 5260 37510
rect 5316 37508 5340 37510
rect 5396 37508 5420 37510
rect 5476 37508 5482 37510
rect 5174 37499 5482 37508
rect 4066 36816 4122 36825
rect 4122 36774 4200 36802
rect 4066 36751 4122 36760
rect 4172 30190 4200 36774
rect 5174 36476 5482 36485
rect 5174 36474 5180 36476
rect 5236 36474 5260 36476
rect 5316 36474 5340 36476
rect 5396 36474 5420 36476
rect 5476 36474 5482 36476
rect 5236 36422 5238 36474
rect 5418 36422 5420 36474
rect 5174 36420 5180 36422
rect 5236 36420 5260 36422
rect 5316 36420 5340 36422
rect 5396 36420 5420 36422
rect 5476 36420 5482 36422
rect 5174 36411 5482 36420
rect 5174 35388 5482 35397
rect 5174 35386 5180 35388
rect 5236 35386 5260 35388
rect 5316 35386 5340 35388
rect 5396 35386 5420 35388
rect 5476 35386 5482 35388
rect 5236 35334 5238 35386
rect 5418 35334 5420 35386
rect 5174 35332 5180 35334
rect 5236 35332 5260 35334
rect 5316 35332 5340 35334
rect 5396 35332 5420 35334
rect 5476 35332 5482 35334
rect 5174 35323 5482 35332
rect 5174 34300 5482 34309
rect 5174 34298 5180 34300
rect 5236 34298 5260 34300
rect 5316 34298 5340 34300
rect 5396 34298 5420 34300
rect 5476 34298 5482 34300
rect 5236 34246 5238 34298
rect 5418 34246 5420 34298
rect 5174 34244 5180 34246
rect 5236 34244 5260 34246
rect 5316 34244 5340 34246
rect 5396 34244 5420 34246
rect 5476 34244 5482 34246
rect 5174 34235 5482 34244
rect 5174 33212 5482 33221
rect 5174 33210 5180 33212
rect 5236 33210 5260 33212
rect 5316 33210 5340 33212
rect 5396 33210 5420 33212
rect 5476 33210 5482 33212
rect 5236 33158 5238 33210
rect 5418 33158 5420 33210
rect 5174 33156 5180 33158
rect 5236 33156 5260 33158
rect 5316 33156 5340 33158
rect 5396 33156 5420 33158
rect 5476 33156 5482 33158
rect 5174 33147 5482 33156
rect 5174 32124 5482 32133
rect 5174 32122 5180 32124
rect 5236 32122 5260 32124
rect 5316 32122 5340 32124
rect 5396 32122 5420 32124
rect 5476 32122 5482 32124
rect 5236 32070 5238 32122
rect 5418 32070 5420 32122
rect 5174 32068 5180 32070
rect 5236 32068 5260 32070
rect 5316 32068 5340 32070
rect 5396 32068 5420 32070
rect 5476 32068 5482 32070
rect 5174 32059 5482 32068
rect 5174 31036 5482 31045
rect 5174 31034 5180 31036
rect 5236 31034 5260 31036
rect 5316 31034 5340 31036
rect 5396 31034 5420 31036
rect 5476 31034 5482 31036
rect 5236 30982 5238 31034
rect 5418 30982 5420 31034
rect 5174 30980 5180 30982
rect 5236 30980 5260 30982
rect 5316 30980 5340 30982
rect 5396 30980 5420 30982
rect 5476 30980 5482 30982
rect 5174 30971 5482 30980
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 5174 29948 5482 29957
rect 5174 29946 5180 29948
rect 5236 29946 5260 29948
rect 5316 29946 5340 29948
rect 5396 29946 5420 29948
rect 5476 29946 5482 29948
rect 5236 29894 5238 29946
rect 5418 29894 5420 29946
rect 5174 29892 5180 29894
rect 5236 29892 5260 29894
rect 5316 29892 5340 29894
rect 5396 29892 5420 29894
rect 5476 29892 5482 29894
rect 5174 29883 5482 29892
rect 5174 28860 5482 28869
rect 5174 28858 5180 28860
rect 5236 28858 5260 28860
rect 5316 28858 5340 28860
rect 5396 28858 5420 28860
rect 5476 28858 5482 28860
rect 5236 28806 5238 28858
rect 5418 28806 5420 28858
rect 5174 28804 5180 28806
rect 5236 28804 5260 28806
rect 5316 28804 5340 28806
rect 5396 28804 5420 28806
rect 5476 28804 5482 28806
rect 5174 28795 5482 28804
rect 5174 27772 5482 27781
rect 5174 27770 5180 27772
rect 5236 27770 5260 27772
rect 5316 27770 5340 27772
rect 5396 27770 5420 27772
rect 5476 27770 5482 27772
rect 5236 27718 5238 27770
rect 5418 27718 5420 27770
rect 5174 27716 5180 27718
rect 5236 27716 5260 27718
rect 5316 27716 5340 27718
rect 5396 27716 5420 27718
rect 5476 27716 5482 27718
rect 5174 27707 5482 27716
rect 5174 26684 5482 26693
rect 5174 26682 5180 26684
rect 5236 26682 5260 26684
rect 5316 26682 5340 26684
rect 5396 26682 5420 26684
rect 5476 26682 5482 26684
rect 5236 26630 5238 26682
rect 5418 26630 5420 26682
rect 5174 26628 5180 26630
rect 5236 26628 5260 26630
rect 5316 26628 5340 26630
rect 5396 26628 5420 26630
rect 5476 26628 5482 26630
rect 5174 26619 5482 26628
rect 3608 25968 3660 25974
rect 3608 25910 3660 25916
rect 5174 25596 5482 25605
rect 5174 25594 5180 25596
rect 5236 25594 5260 25596
rect 5316 25594 5340 25596
rect 5396 25594 5420 25596
rect 5476 25594 5482 25596
rect 5236 25542 5238 25594
rect 5418 25542 5420 25594
rect 5174 25540 5180 25542
rect 5236 25540 5260 25542
rect 5316 25540 5340 25542
rect 5396 25540 5420 25542
rect 5476 25540 5482 25542
rect 5174 25531 5482 25540
rect 5174 24508 5482 24517
rect 5174 24506 5180 24508
rect 5236 24506 5260 24508
rect 5316 24506 5340 24508
rect 5396 24506 5420 24508
rect 5476 24506 5482 24508
rect 5236 24454 5238 24506
rect 5418 24454 5420 24506
rect 5174 24452 5180 24454
rect 5236 24452 5260 24454
rect 5316 24452 5340 24454
rect 5396 24452 5420 24454
rect 5476 24452 5482 24454
rect 5174 24443 5482 24452
rect 5174 23420 5482 23429
rect 5174 23418 5180 23420
rect 5236 23418 5260 23420
rect 5316 23418 5340 23420
rect 5396 23418 5420 23420
rect 5476 23418 5482 23420
rect 5236 23366 5238 23418
rect 5418 23366 5420 23418
rect 5174 23364 5180 23366
rect 5236 23364 5260 23366
rect 5316 23364 5340 23366
rect 5396 23364 5420 23366
rect 5476 23364 5482 23366
rect 5174 23355 5482 23364
rect 5174 22332 5482 22341
rect 5174 22330 5180 22332
rect 5236 22330 5260 22332
rect 5316 22330 5340 22332
rect 5396 22330 5420 22332
rect 5476 22330 5482 22332
rect 5236 22278 5238 22330
rect 5418 22278 5420 22330
rect 5174 22276 5180 22278
rect 5236 22276 5260 22278
rect 5316 22276 5340 22278
rect 5396 22276 5420 22278
rect 5476 22276 5482 22278
rect 5174 22267 5482 22276
rect 5174 21244 5482 21253
rect 5174 21242 5180 21244
rect 5236 21242 5260 21244
rect 5316 21242 5340 21244
rect 5396 21242 5420 21244
rect 5476 21242 5482 21244
rect 5236 21190 5238 21242
rect 5418 21190 5420 21242
rect 5174 21188 5180 21190
rect 5236 21188 5260 21190
rect 5316 21188 5340 21190
rect 5396 21188 5420 21190
rect 5476 21188 5482 21190
rect 5174 21179 5482 21188
rect 5174 20156 5482 20165
rect 5174 20154 5180 20156
rect 5236 20154 5260 20156
rect 5316 20154 5340 20156
rect 5396 20154 5420 20156
rect 5476 20154 5482 20156
rect 5236 20102 5238 20154
rect 5418 20102 5420 20154
rect 5174 20100 5180 20102
rect 5236 20100 5260 20102
rect 5316 20100 5340 20102
rect 5396 20100 5420 20102
rect 5476 20100 5482 20102
rect 5174 20091 5482 20100
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 6276 19168 6328 19174
rect 3422 19136 3478 19145
rect 6276 19110 6328 19116
rect 3422 19071 3478 19080
rect 3436 18630 3464 19071
rect 5174 19068 5482 19077
rect 5174 19066 5180 19068
rect 5236 19066 5260 19068
rect 5316 19066 5340 19068
rect 5396 19066 5420 19068
rect 5476 19066 5482 19068
rect 5236 19014 5238 19066
rect 5418 19014 5420 19066
rect 5174 19012 5180 19014
rect 5236 19012 5260 19014
rect 5316 19012 5340 19014
rect 5396 19012 5420 19014
rect 5476 19012 5482 19014
rect 5174 19003 5482 19012
rect 6288 18834 6316 19110
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3422 18456 3478 18465
rect 3422 18391 3478 18400
rect 3436 18222 3464 18391
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 5092 17746 5120 18702
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18426 6684 18634
rect 6748 18426 6776 37810
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 5174 17980 5482 17989
rect 5174 17978 5180 17980
rect 5236 17978 5260 17980
rect 5316 17978 5340 17980
rect 5396 17978 5420 17980
rect 5476 17978 5482 17980
rect 5236 17926 5238 17978
rect 5418 17926 5420 17978
rect 5174 17924 5180 17926
rect 5236 17924 5260 17926
rect 5316 17924 5340 17926
rect 5396 17924 5420 17926
rect 5476 17924 5482 17926
rect 5174 17915 5482 17924
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5368 17338 5396 17546
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 3332 17128 3384 17134
rect 3238 17096 3294 17105
rect 3332 17070 3384 17076
rect 3238 17031 3294 17040
rect 3252 16590 3280 17031
rect 5174 16892 5482 16901
rect 5174 16890 5180 16892
rect 5236 16890 5260 16892
rect 5316 16890 5340 16892
rect 5396 16890 5420 16892
rect 5476 16890 5482 16892
rect 5236 16838 5238 16890
rect 5418 16838 5420 16890
rect 5174 16836 5180 16838
rect 5236 16836 5260 16838
rect 5316 16836 5340 16838
rect 5396 16836 5420 16838
rect 5476 16836 5482 16838
rect 5174 16827 5482 16836
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4066 15736 4122 15745
rect 4066 15671 4122 15680
rect 4080 15638 4108 15671
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4264 15570 4292 15846
rect 5174 15804 5482 15813
rect 5174 15802 5180 15804
rect 5236 15802 5260 15804
rect 5316 15802 5340 15804
rect 5396 15802 5420 15804
rect 5476 15802 5482 15804
rect 5236 15750 5238 15802
rect 5418 15750 5420 15802
rect 5174 15748 5180 15750
rect 5236 15748 5260 15750
rect 5316 15748 5340 15750
rect 5396 15748 5420 15750
rect 5476 15748 5482 15750
rect 5174 15739 5482 15748
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4436 15428 4488 15434
rect 4436 15370 4488 15376
rect 4448 15162 4476 15370
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5174 14716 5482 14725
rect 5174 14714 5180 14716
rect 5236 14714 5260 14716
rect 5316 14714 5340 14716
rect 5396 14714 5420 14716
rect 5476 14714 5482 14716
rect 5236 14662 5238 14714
rect 5418 14662 5420 14714
rect 5174 14660 5180 14662
rect 5236 14660 5260 14662
rect 5316 14660 5340 14662
rect 5396 14660 5420 14662
rect 5476 14660 5482 14662
rect 5174 14651 5482 14660
rect 5174 13628 5482 13637
rect 5174 13626 5180 13628
rect 5236 13626 5260 13628
rect 5316 13626 5340 13628
rect 5396 13626 5420 13628
rect 5476 13626 5482 13628
rect 5236 13574 5238 13626
rect 5418 13574 5420 13626
rect 5174 13572 5180 13574
rect 5236 13572 5260 13574
rect 5316 13572 5340 13574
rect 5396 13572 5420 13574
rect 5476 13572 5482 13574
rect 5174 13563 5482 13572
rect 5644 12986 5672 14962
rect 6564 13938 6592 18022
rect 6840 17746 6868 38542
rect 7116 37874 7144 41200
rect 7104 37868 7156 37874
rect 7104 37810 7156 37816
rect 7300 26234 7328 41262
rect 7576 41154 7604 41262
rect 7718 41200 7830 42000
rect 8362 41200 8474 42000
rect 9006 41200 9118 42000
rect 9650 41200 9762 42000
rect 10938 41200 11050 42000
rect 11582 41200 11694 42000
rect 12226 41200 12338 42000
rect 12870 41200 12982 42000
rect 13514 41200 13626 42000
rect 14158 41200 14270 42000
rect 14802 41200 14914 42000
rect 15446 41200 15558 42000
rect 16090 41200 16202 42000
rect 17378 41200 17490 42000
rect 18022 41200 18134 42000
rect 18666 41200 18778 42000
rect 19310 41200 19422 42000
rect 19954 41200 20066 42000
rect 20180 41262 20484 41290
rect 7760 41154 7788 41200
rect 7576 41126 7788 41154
rect 7840 39432 7892 39438
rect 7840 39374 7892 39380
rect 7852 38962 7880 39374
rect 7840 38956 7892 38962
rect 7840 38898 7892 38904
rect 8404 38894 8432 41200
rect 8024 38888 8076 38894
rect 8024 38830 8076 38836
rect 8392 38888 8444 38894
rect 8392 38830 8444 38836
rect 8036 38554 8064 38830
rect 8024 38548 8076 38554
rect 8024 38490 8076 38496
rect 9048 38486 9076 41200
rect 13622 39740 13930 39749
rect 13622 39738 13628 39740
rect 13684 39738 13708 39740
rect 13764 39738 13788 39740
rect 13844 39738 13868 39740
rect 13924 39738 13930 39740
rect 13684 39686 13686 39738
rect 13866 39686 13868 39738
rect 13622 39684 13628 39686
rect 13684 39684 13708 39686
rect 13764 39684 13788 39686
rect 13844 39684 13868 39686
rect 13924 39684 13930 39686
rect 13622 39675 13930 39684
rect 9398 39196 9706 39205
rect 9398 39194 9404 39196
rect 9460 39194 9484 39196
rect 9540 39194 9564 39196
rect 9620 39194 9644 39196
rect 9700 39194 9706 39196
rect 9460 39142 9462 39194
rect 9642 39142 9644 39194
rect 9398 39140 9404 39142
rect 9460 39140 9484 39142
rect 9540 39140 9564 39142
rect 9620 39140 9644 39142
rect 9700 39140 9706 39142
rect 9398 39131 9706 39140
rect 13622 38652 13930 38661
rect 13622 38650 13628 38652
rect 13684 38650 13708 38652
rect 13764 38650 13788 38652
rect 13844 38650 13868 38652
rect 13924 38650 13930 38652
rect 13684 38598 13686 38650
rect 13866 38598 13868 38650
rect 13622 38596 13628 38598
rect 13684 38596 13708 38598
rect 13764 38596 13788 38598
rect 13844 38596 13868 38598
rect 13924 38596 13930 38598
rect 13622 38587 13930 38596
rect 9036 38480 9088 38486
rect 9036 38422 9088 38428
rect 9398 38108 9706 38117
rect 9398 38106 9404 38108
rect 9460 38106 9484 38108
rect 9540 38106 9564 38108
rect 9620 38106 9644 38108
rect 9700 38106 9706 38108
rect 9460 38054 9462 38106
rect 9642 38054 9644 38106
rect 9398 38052 9404 38054
rect 9460 38052 9484 38054
rect 9540 38052 9564 38054
rect 9620 38052 9644 38054
rect 9700 38052 9706 38054
rect 9398 38043 9706 38052
rect 10416 37868 10468 37874
rect 10416 37810 10468 37816
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8404 37262 8432 37606
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 7380 37188 7432 37194
rect 7380 37130 7432 37136
rect 7392 36922 7420 37130
rect 9398 37020 9706 37029
rect 9398 37018 9404 37020
rect 9460 37018 9484 37020
rect 9540 37018 9564 37020
rect 9620 37018 9644 37020
rect 9700 37018 9706 37020
rect 9460 36966 9462 37018
rect 9642 36966 9644 37018
rect 9398 36964 9404 36966
rect 9460 36964 9484 36966
rect 9540 36964 9564 36966
rect 9620 36964 9644 36966
rect 9700 36964 9706 36966
rect 9398 36955 9706 36964
rect 7380 36916 7432 36922
rect 7380 36858 7432 36864
rect 9398 35932 9706 35941
rect 9398 35930 9404 35932
rect 9460 35930 9484 35932
rect 9540 35930 9564 35932
rect 9620 35930 9644 35932
rect 9700 35930 9706 35932
rect 9460 35878 9462 35930
rect 9642 35878 9644 35930
rect 9398 35876 9404 35878
rect 9460 35876 9484 35878
rect 9540 35876 9564 35878
rect 9620 35876 9644 35878
rect 9700 35876 9706 35878
rect 9398 35867 9706 35876
rect 9398 34844 9706 34853
rect 9398 34842 9404 34844
rect 9460 34842 9484 34844
rect 9540 34842 9564 34844
rect 9620 34842 9644 34844
rect 9700 34842 9706 34844
rect 9460 34790 9462 34842
rect 9642 34790 9644 34842
rect 9398 34788 9404 34790
rect 9460 34788 9484 34790
rect 9540 34788 9564 34790
rect 9620 34788 9644 34790
rect 9700 34788 9706 34790
rect 9398 34779 9706 34788
rect 9864 34400 9916 34406
rect 9864 34342 9916 34348
rect 9876 34066 9904 34342
rect 9864 34060 9916 34066
rect 9864 34002 9916 34008
rect 10232 33924 10284 33930
rect 10232 33866 10284 33872
rect 9398 33756 9706 33765
rect 9398 33754 9404 33756
rect 9460 33754 9484 33756
rect 9540 33754 9564 33756
rect 9620 33754 9644 33756
rect 9700 33754 9706 33756
rect 9460 33702 9462 33754
rect 9642 33702 9644 33754
rect 9398 33700 9404 33702
rect 9460 33700 9484 33702
rect 9540 33700 9564 33702
rect 9620 33700 9644 33702
rect 9700 33700 9706 33702
rect 9398 33691 9706 33700
rect 10244 33658 10272 33866
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10324 33516 10376 33522
rect 10324 33458 10376 33464
rect 9398 32668 9706 32677
rect 9398 32666 9404 32668
rect 9460 32666 9484 32668
rect 9540 32666 9564 32668
rect 9620 32666 9644 32668
rect 9700 32666 9706 32668
rect 9460 32614 9462 32666
rect 9642 32614 9644 32666
rect 9398 32612 9404 32614
rect 9460 32612 9484 32614
rect 9540 32612 9564 32614
rect 9620 32612 9644 32614
rect 9700 32612 9706 32614
rect 9398 32603 9706 32612
rect 9398 31580 9706 31589
rect 9398 31578 9404 31580
rect 9460 31578 9484 31580
rect 9540 31578 9564 31580
rect 9620 31578 9644 31580
rect 9700 31578 9706 31580
rect 9460 31526 9462 31578
rect 9642 31526 9644 31578
rect 9398 31524 9404 31526
rect 9460 31524 9484 31526
rect 9540 31524 9564 31526
rect 9620 31524 9644 31526
rect 9700 31524 9706 31526
rect 9398 31515 9706 31524
rect 9398 30492 9706 30501
rect 9398 30490 9404 30492
rect 9460 30490 9484 30492
rect 9540 30490 9564 30492
rect 9620 30490 9644 30492
rect 9700 30490 9706 30492
rect 9460 30438 9462 30490
rect 9642 30438 9644 30490
rect 9398 30436 9404 30438
rect 9460 30436 9484 30438
rect 9540 30436 9564 30438
rect 9620 30436 9644 30438
rect 9700 30436 9706 30438
rect 9398 30427 9706 30436
rect 9398 29404 9706 29413
rect 9398 29402 9404 29404
rect 9460 29402 9484 29404
rect 9540 29402 9564 29404
rect 9620 29402 9644 29404
rect 9700 29402 9706 29404
rect 9460 29350 9462 29402
rect 9642 29350 9644 29402
rect 9398 29348 9404 29350
rect 9460 29348 9484 29350
rect 9540 29348 9564 29350
rect 9620 29348 9644 29350
rect 9700 29348 9706 29350
rect 9398 29339 9706 29348
rect 9398 28316 9706 28325
rect 9398 28314 9404 28316
rect 9460 28314 9484 28316
rect 9540 28314 9564 28316
rect 9620 28314 9644 28316
rect 9700 28314 9706 28316
rect 9460 28262 9462 28314
rect 9642 28262 9644 28314
rect 9398 28260 9404 28262
rect 9460 28260 9484 28262
rect 9540 28260 9564 28262
rect 9620 28260 9644 28262
rect 9700 28260 9706 28262
rect 9398 28251 9706 28260
rect 9398 27228 9706 27237
rect 9398 27226 9404 27228
rect 9460 27226 9484 27228
rect 9540 27226 9564 27228
rect 9620 27226 9644 27228
rect 9700 27226 9706 27228
rect 9460 27174 9462 27226
rect 9642 27174 9644 27226
rect 9398 27172 9404 27174
rect 9460 27172 9484 27174
rect 9540 27172 9564 27174
rect 9620 27172 9644 27174
rect 9700 27172 9706 27174
rect 9398 27163 9706 27172
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 6932 26206 7328 26234
rect 6932 17814 6960 26206
rect 8864 25974 8892 26318
rect 9398 26140 9706 26149
rect 9398 26138 9404 26140
rect 9460 26138 9484 26140
rect 9540 26138 9564 26140
rect 9620 26138 9644 26140
rect 9700 26138 9706 26140
rect 9460 26086 9462 26138
rect 9642 26086 9644 26138
rect 9398 26084 9404 26086
rect 9460 26084 9484 26086
rect 9540 26084 9564 26086
rect 9620 26084 9644 26086
rect 9700 26084 9706 26086
rect 9398 26075 9706 26084
rect 8852 25968 8904 25974
rect 8852 25910 8904 25916
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 9048 25498 9076 25774
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9968 25362 9996 25638
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 7668 24818 7696 25230
rect 8392 24948 8444 24954
rect 8392 24890 8444 24896
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 8404 24750 8432 24890
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8312 24410 8340 24686
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8496 19378 8524 20198
rect 8680 19446 8708 20198
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 7852 17542 7880 18226
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6196 13462 6224 13806
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5644 12850 5672 12922
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4066 11656 4122 11665
rect 4172 11642 4200 12718
rect 5174 12540 5482 12549
rect 5174 12538 5180 12540
rect 5236 12538 5260 12540
rect 5316 12538 5340 12540
rect 5396 12538 5420 12540
rect 5476 12538 5482 12540
rect 5236 12486 5238 12538
rect 5418 12486 5420 12538
rect 5174 12484 5180 12486
rect 5236 12484 5260 12486
rect 5316 12484 5340 12486
rect 5396 12484 5420 12486
rect 5476 12484 5482 12486
rect 5174 12475 5482 12484
rect 4122 11614 4200 11642
rect 4066 11591 4122 11600
rect 5174 11452 5482 11461
rect 5174 11450 5180 11452
rect 5236 11450 5260 11452
rect 5316 11450 5340 11452
rect 5396 11450 5420 11452
rect 5476 11450 5482 11452
rect 5236 11398 5238 11450
rect 5418 11398 5420 11450
rect 5174 11396 5180 11398
rect 5236 11396 5260 11398
rect 5316 11396 5340 11398
rect 5396 11396 5420 11398
rect 5476 11396 5482 11398
rect 5174 11387 5482 11396
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3148 8288 3200 8294
rect 3146 8256 3148 8265
rect 3200 8256 3202 8265
rect 3146 8191 3202 8200
rect 3146 7576 3202 7585
rect 3146 7511 3202 7520
rect 3160 7342 3188 7511
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2792 3058 2820 3470
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2608 800 2636 2858
rect 2976 2650 3004 2926
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2446 3096 6734
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3252 800 3280 3334
rect 3344 1465 3372 11018
rect 5174 10364 5482 10373
rect 5174 10362 5180 10364
rect 5236 10362 5260 10364
rect 5316 10362 5340 10364
rect 5396 10362 5420 10364
rect 5476 10362 5482 10364
rect 5236 10310 5238 10362
rect 5418 10310 5420 10362
rect 5174 10308 5180 10310
rect 5236 10308 5260 10310
rect 5316 10308 5340 10310
rect 5396 10308 5420 10310
rect 5476 10308 5482 10310
rect 5174 10299 5482 10308
rect 5174 9276 5482 9285
rect 5174 9274 5180 9276
rect 5236 9274 5260 9276
rect 5316 9274 5340 9276
rect 5396 9274 5420 9276
rect 5476 9274 5482 9276
rect 5236 9222 5238 9274
rect 5418 9222 5420 9274
rect 5174 9220 5180 9222
rect 5236 9220 5260 9222
rect 5316 9220 5340 9222
rect 5396 9220 5420 9222
rect 5476 9220 5482 9222
rect 5174 9211 5482 9220
rect 5174 8188 5482 8197
rect 5174 8186 5180 8188
rect 5236 8186 5260 8188
rect 5316 8186 5340 8188
rect 5396 8186 5420 8188
rect 5476 8186 5482 8188
rect 5236 8134 5238 8186
rect 5418 8134 5420 8186
rect 5174 8132 5180 8134
rect 5236 8132 5260 8134
rect 5316 8132 5340 8134
rect 5396 8132 5420 8134
rect 5476 8132 5482 8134
rect 5174 8123 5482 8132
rect 6564 7410 6592 13874
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13258 6960 13806
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10810 7144 11018
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7300 10606 7328 11086
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 5174 7100 5482 7109
rect 5174 7098 5180 7100
rect 5236 7098 5260 7100
rect 5316 7098 5340 7100
rect 5396 7098 5420 7100
rect 5476 7098 5482 7100
rect 5236 7046 5238 7098
rect 5418 7046 5420 7098
rect 5174 7044 5180 7046
rect 5236 7044 5260 7046
rect 5316 7044 5340 7046
rect 5396 7044 5420 7046
rect 5476 7044 5482 7046
rect 5174 7035 5482 7044
rect 6564 6914 6592 7346
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6564 6886 6684 6914
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5174 6012 5482 6021
rect 5174 6010 5180 6012
rect 5236 6010 5260 6012
rect 5316 6010 5340 6012
rect 5396 6010 5420 6012
rect 5476 6010 5482 6012
rect 5236 5958 5238 6010
rect 5418 5958 5420 6010
rect 5174 5956 5180 5958
rect 5236 5956 5260 5958
rect 5316 5956 5340 5958
rect 5396 5956 5420 5958
rect 5476 5956 5482 5958
rect 5174 5947 5482 5956
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3436 5302 3464 5471
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 5174 4924 5482 4933
rect 5174 4922 5180 4924
rect 5236 4922 5260 4924
rect 5316 4922 5340 4924
rect 5396 4922 5420 4924
rect 5476 4922 5482 4924
rect 5236 4870 5238 4922
rect 5418 4870 5420 4922
rect 5174 4868 5180 4870
rect 5236 4868 5260 4870
rect 5316 4868 5340 4870
rect 5396 4868 5420 4870
rect 5476 4868 5482 4870
rect 5174 4859 5482 4868
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3436 4185 3464 4694
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 3505 3464 4014
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3422 3496 3478 3505
rect 3422 3431 3478 3440
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3436 2825 3464 2858
rect 3422 2816 3478 2825
rect 3422 2751 3478 2760
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 2145 3464 2246
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3896 800 3924 3946
rect 5174 3836 5482 3845
rect 5174 3834 5180 3836
rect 5236 3834 5260 3836
rect 5316 3834 5340 3836
rect 5396 3834 5420 3836
rect 5476 3834 5482 3836
rect 5236 3782 5238 3834
rect 5418 3782 5420 3834
rect 5174 3780 5180 3782
rect 5236 3780 5260 3782
rect 5316 3780 5340 3782
rect 5396 3780 5420 3782
rect 5476 3780 5482 3782
rect 5174 3771 5482 3780
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 800 4568 2790
rect 5092 1850 5120 3538
rect 5552 2854 5580 4490
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5174 2748 5482 2757
rect 5174 2746 5180 2748
rect 5236 2746 5260 2748
rect 5316 2746 5340 2748
rect 5396 2746 5420 2748
rect 5476 2746 5482 2748
rect 5236 2694 5238 2746
rect 5418 2694 5420 2746
rect 5174 2692 5180 2694
rect 5236 2692 5260 2694
rect 5316 2692 5340 2694
rect 5396 2692 5420 2694
rect 5476 2692 5482 2694
rect 5174 2683 5482 2692
rect 5644 2310 5672 6122
rect 6196 3398 6224 6666
rect 6656 4690 6684 6886
rect 7116 6730 7144 7142
rect 7300 6866 7328 7142
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7116 5234 7144 5714
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 7116 4146 7144 4966
rect 7392 4622 7420 17478
rect 8128 6914 8156 18634
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18154 9076 18566
rect 9140 18290 9168 19790
rect 9324 18970 9352 25230
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 9398 25052 9706 25061
rect 9398 25050 9404 25052
rect 9460 25050 9484 25052
rect 9540 25050 9564 25052
rect 9620 25050 9644 25052
rect 9700 25050 9706 25052
rect 9460 24998 9462 25050
rect 9642 24998 9644 25050
rect 9398 24996 9404 24998
rect 9460 24996 9484 24998
rect 9540 24996 9564 24998
rect 9620 24996 9644 24998
rect 9700 24996 9706 24998
rect 9398 24987 9706 24996
rect 10152 24954 10180 25162
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 9398 23964 9706 23973
rect 9398 23962 9404 23964
rect 9460 23962 9484 23964
rect 9540 23962 9564 23964
rect 9620 23962 9644 23964
rect 9700 23962 9706 23964
rect 9460 23910 9462 23962
rect 9642 23910 9644 23962
rect 9398 23908 9404 23910
rect 9460 23908 9484 23910
rect 9540 23908 9564 23910
rect 9620 23908 9644 23910
rect 9700 23908 9706 23910
rect 9398 23899 9706 23908
rect 9398 22876 9706 22885
rect 9398 22874 9404 22876
rect 9460 22874 9484 22876
rect 9540 22874 9564 22876
rect 9620 22874 9644 22876
rect 9700 22874 9706 22876
rect 9460 22822 9462 22874
rect 9642 22822 9644 22874
rect 9398 22820 9404 22822
rect 9460 22820 9484 22822
rect 9540 22820 9564 22822
rect 9620 22820 9644 22822
rect 9700 22820 9706 22822
rect 9398 22811 9706 22820
rect 9398 21788 9706 21797
rect 9398 21786 9404 21788
rect 9460 21786 9484 21788
rect 9540 21786 9564 21788
rect 9620 21786 9644 21788
rect 9700 21786 9706 21788
rect 9460 21734 9462 21786
rect 9642 21734 9644 21786
rect 9398 21732 9404 21734
rect 9460 21732 9484 21734
rect 9540 21732 9564 21734
rect 9620 21732 9644 21734
rect 9700 21732 9706 21734
rect 9398 21723 9706 21732
rect 9398 20700 9706 20709
rect 9398 20698 9404 20700
rect 9460 20698 9484 20700
rect 9540 20698 9564 20700
rect 9620 20698 9644 20700
rect 9700 20698 9706 20700
rect 9460 20646 9462 20698
rect 9642 20646 9644 20698
rect 9398 20644 9404 20646
rect 9460 20644 9484 20646
rect 9540 20644 9564 20646
rect 9620 20644 9644 20646
rect 9700 20644 9706 20646
rect 9398 20635 9706 20644
rect 10336 20534 10364 33458
rect 10428 25362 10456 37810
rect 13622 37564 13930 37573
rect 13622 37562 13628 37564
rect 13684 37562 13708 37564
rect 13764 37562 13788 37564
rect 13844 37562 13868 37564
rect 13924 37562 13930 37564
rect 13684 37510 13686 37562
rect 13866 37510 13868 37562
rect 13622 37508 13628 37510
rect 13684 37508 13708 37510
rect 13764 37508 13788 37510
rect 13844 37508 13868 37510
rect 13924 37508 13930 37510
rect 13622 37499 13930 37508
rect 13622 36476 13930 36485
rect 13622 36474 13628 36476
rect 13684 36474 13708 36476
rect 13764 36474 13788 36476
rect 13844 36474 13868 36476
rect 13924 36474 13930 36476
rect 13684 36422 13686 36474
rect 13866 36422 13868 36474
rect 13622 36420 13628 36422
rect 13684 36420 13708 36422
rect 13764 36420 13788 36422
rect 13844 36420 13868 36422
rect 13924 36420 13930 36422
rect 13622 36411 13930 36420
rect 13622 35388 13930 35397
rect 13622 35386 13628 35388
rect 13684 35386 13708 35388
rect 13764 35386 13788 35388
rect 13844 35386 13868 35388
rect 13924 35386 13930 35388
rect 13684 35334 13686 35386
rect 13866 35334 13868 35386
rect 13622 35332 13628 35334
rect 13684 35332 13708 35334
rect 13764 35332 13788 35334
rect 13844 35332 13868 35334
rect 13924 35332 13930 35334
rect 13622 35323 13930 35332
rect 13622 34300 13930 34309
rect 13622 34298 13628 34300
rect 13684 34298 13708 34300
rect 13764 34298 13788 34300
rect 13844 34298 13868 34300
rect 13924 34298 13930 34300
rect 13684 34246 13686 34298
rect 13866 34246 13868 34298
rect 13622 34244 13628 34246
rect 13684 34244 13708 34246
rect 13764 34244 13788 34246
rect 13844 34244 13868 34246
rect 13924 34244 13930 34246
rect 13622 34235 13930 34244
rect 13622 33212 13930 33221
rect 13622 33210 13628 33212
rect 13684 33210 13708 33212
rect 13764 33210 13788 33212
rect 13844 33210 13868 33212
rect 13924 33210 13930 33212
rect 13684 33158 13686 33210
rect 13866 33158 13868 33210
rect 13622 33156 13628 33158
rect 13684 33156 13708 33158
rect 13764 33156 13788 33158
rect 13844 33156 13868 33158
rect 13924 33156 13930 33158
rect 13622 33147 13930 33156
rect 13622 32124 13930 32133
rect 13622 32122 13628 32124
rect 13684 32122 13708 32124
rect 13764 32122 13788 32124
rect 13844 32122 13868 32124
rect 13924 32122 13930 32124
rect 13684 32070 13686 32122
rect 13866 32070 13868 32122
rect 13622 32068 13628 32070
rect 13684 32068 13708 32070
rect 13764 32068 13788 32070
rect 13844 32068 13868 32070
rect 13924 32068 13930 32070
rect 13622 32059 13930 32068
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10980 30122 11008 31758
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11716 30938 11744 31214
rect 13622 31036 13930 31045
rect 13622 31034 13628 31036
rect 13684 31034 13708 31036
rect 13764 31034 13788 31036
rect 13844 31034 13868 31036
rect 13924 31034 13930 31036
rect 13684 30982 13686 31034
rect 13866 30982 13868 31034
rect 13622 30980 13628 30982
rect 13684 30980 13708 30982
rect 13764 30980 13788 30982
rect 13844 30980 13868 30982
rect 13924 30980 13930 30982
rect 13622 30971 13930 30980
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 11808 30258 11836 30670
rect 14292 30258 14320 30670
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14844 30190 14872 41200
rect 16132 39522 16160 41200
rect 16132 39494 16252 39522
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 16132 38418 16160 39374
rect 16120 38412 16172 38418
rect 16120 38354 16172 38360
rect 16224 38214 16252 39494
rect 17040 39432 17092 39438
rect 17040 39374 17092 39380
rect 16948 39364 17000 39370
rect 16948 39306 17000 39312
rect 16960 38962 16988 39306
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 17052 38826 17080 39374
rect 17132 39296 17184 39302
rect 17132 39238 17184 39244
rect 17144 39030 17172 39238
rect 17132 39024 17184 39030
rect 17132 38966 17184 38972
rect 17420 38894 17448 41200
rect 18064 39302 18092 41200
rect 18052 39296 18104 39302
rect 18052 39238 18104 39244
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 17846 39196 18154 39205
rect 17846 39194 17852 39196
rect 17908 39194 17932 39196
rect 17988 39194 18012 39196
rect 18068 39194 18092 39196
rect 18148 39194 18154 39196
rect 17908 39142 17910 39194
rect 18090 39142 18092 39194
rect 17846 39140 17852 39142
rect 17908 39140 17932 39142
rect 17988 39140 18012 39142
rect 18068 39140 18092 39142
rect 18148 39140 18154 39142
rect 17846 39131 18154 39140
rect 17408 38888 17460 38894
rect 17408 38830 17460 38836
rect 17040 38820 17092 38826
rect 17040 38762 17092 38768
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16592 38418 16620 38694
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16856 38412 16908 38418
rect 16856 38354 16908 38360
rect 16868 38214 16896 38354
rect 16212 38208 16264 38214
rect 16212 38150 16264 38156
rect 16856 38208 16908 38214
rect 16856 38150 16908 38156
rect 17052 32978 17080 38762
rect 17846 38108 18154 38117
rect 17846 38106 17852 38108
rect 17908 38106 17932 38108
rect 17988 38106 18012 38108
rect 18068 38106 18092 38108
rect 18148 38106 18154 38108
rect 17908 38054 17910 38106
rect 18090 38054 18092 38106
rect 17846 38052 17852 38054
rect 17908 38052 17932 38054
rect 17988 38052 18012 38054
rect 18068 38052 18092 38054
rect 18148 38052 18154 38054
rect 17846 38043 18154 38052
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 17846 37020 18154 37029
rect 17846 37018 17852 37020
rect 17908 37018 17932 37020
rect 17988 37018 18012 37020
rect 18068 37018 18092 37020
rect 18148 37018 18154 37020
rect 17908 36966 17910 37018
rect 18090 36966 18092 37018
rect 17846 36964 17852 36966
rect 17908 36964 17932 36966
rect 17988 36964 18012 36966
rect 18068 36964 18092 36966
rect 18148 36964 18154 36966
rect 17846 36955 18154 36964
rect 18432 36786 18460 37198
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 17316 36576 17368 36582
rect 17316 36518 17368 36524
rect 17328 35698 17356 36518
rect 17512 36174 17540 36722
rect 17500 36168 17552 36174
rect 17500 36110 17552 36116
rect 17316 35692 17368 35698
rect 17316 35634 17368 35640
rect 17040 32972 17092 32978
rect 17040 32914 17092 32920
rect 17052 31890 17080 32914
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 12176 29850 12204 30126
rect 13622 29948 13930 29957
rect 13622 29946 13628 29948
rect 13684 29946 13708 29948
rect 13764 29946 13788 29948
rect 13844 29946 13868 29948
rect 13924 29946 13930 29948
rect 13684 29894 13686 29946
rect 13866 29894 13868 29946
rect 13622 29892 13628 29894
rect 13684 29892 13708 29894
rect 13764 29892 13788 29894
rect 13844 29892 13868 29894
rect 13924 29892 13930 29894
rect 13622 29883 13930 29892
rect 14476 29850 14504 30126
rect 12164 29844 12216 29850
rect 12164 29786 12216 29792
rect 14464 29844 14516 29850
rect 14464 29786 14516 29792
rect 16316 29646 16344 31758
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 13622 28860 13930 28869
rect 13622 28858 13628 28860
rect 13684 28858 13708 28860
rect 13764 28858 13788 28860
rect 13844 28858 13868 28860
rect 13924 28858 13930 28860
rect 13684 28806 13686 28858
rect 13866 28806 13868 28858
rect 13622 28804 13628 28806
rect 13684 28804 13708 28806
rect 13764 28804 13788 28806
rect 13844 28804 13868 28806
rect 13924 28804 13930 28806
rect 13622 28795 13930 28804
rect 13622 27772 13930 27781
rect 13622 27770 13628 27772
rect 13684 27770 13708 27772
rect 13764 27770 13788 27772
rect 13844 27770 13868 27772
rect 13924 27770 13930 27772
rect 13684 27718 13686 27770
rect 13866 27718 13868 27770
rect 13622 27716 13628 27718
rect 13684 27716 13708 27718
rect 13764 27716 13788 27718
rect 13844 27716 13868 27718
rect 13924 27716 13930 27718
rect 13622 27707 13930 27716
rect 13622 26684 13930 26693
rect 13622 26682 13628 26684
rect 13684 26682 13708 26684
rect 13764 26682 13788 26684
rect 13844 26682 13868 26684
rect 13924 26682 13930 26684
rect 13684 26630 13686 26682
rect 13866 26630 13868 26682
rect 13622 26628 13628 26630
rect 13684 26628 13708 26630
rect 13764 26628 13788 26630
rect 13844 26628 13868 26630
rect 13924 26628 13930 26630
rect 13622 26619 13930 26628
rect 13622 25596 13930 25605
rect 13622 25594 13628 25596
rect 13684 25594 13708 25596
rect 13764 25594 13788 25596
rect 13844 25594 13868 25596
rect 13924 25594 13930 25596
rect 13684 25542 13686 25594
rect 13866 25542 13868 25594
rect 13622 25540 13628 25542
rect 13684 25540 13708 25542
rect 13764 25540 13788 25542
rect 13844 25540 13868 25542
rect 13924 25540 13930 25542
rect 13622 25531 13930 25540
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 11072 24206 11100 24754
rect 13622 24508 13930 24517
rect 13622 24506 13628 24508
rect 13684 24506 13708 24508
rect 13764 24506 13788 24508
rect 13844 24506 13868 24508
rect 13924 24506 13930 24508
rect 13684 24454 13686 24506
rect 13866 24454 13868 24506
rect 13622 24452 13628 24454
rect 13684 24452 13708 24454
rect 13764 24452 13788 24454
rect 13844 24452 13868 24454
rect 13924 24452 13930 24454
rect 13622 24443 13930 24452
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 9398 19612 9706 19621
rect 9398 19610 9404 19612
rect 9460 19610 9484 19612
rect 9540 19610 9564 19612
rect 9620 19610 9644 19612
rect 9700 19610 9706 19612
rect 9460 19558 9462 19610
rect 9642 19558 9644 19610
rect 9398 19556 9404 19558
rect 9460 19556 9484 19558
rect 9540 19556 9564 19558
rect 9620 19556 9644 19558
rect 9700 19556 9706 19558
rect 9398 19547 9706 19556
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9324 18766 9352 18906
rect 10244 18834 10272 19110
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9398 18524 9706 18533
rect 9398 18522 9404 18524
rect 9460 18522 9484 18524
rect 9540 18522 9564 18524
rect 9620 18522 9644 18524
rect 9700 18522 9706 18524
rect 9460 18470 9462 18522
rect 9642 18470 9644 18522
rect 9398 18468 9404 18470
rect 9460 18468 9484 18470
rect 9540 18468 9564 18470
rect 9620 18468 9644 18470
rect 9700 18468 9706 18470
rect 9398 18459 9706 18468
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8496 17610 8524 18022
rect 8680 17746 8708 18022
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 9398 17436 9706 17445
rect 9398 17434 9404 17436
rect 9460 17434 9484 17436
rect 9540 17434 9564 17436
rect 9620 17434 9644 17436
rect 9700 17434 9706 17436
rect 9460 17382 9462 17434
rect 9642 17382 9644 17434
rect 9398 17380 9404 17382
rect 9460 17380 9484 17382
rect 9540 17380 9564 17382
rect 9620 17380 9644 17382
rect 9700 17380 9706 17382
rect 9398 17371 9706 17380
rect 9398 16348 9706 16357
rect 9398 16346 9404 16348
rect 9460 16346 9484 16348
rect 9540 16346 9564 16348
rect 9620 16346 9644 16348
rect 9700 16346 9706 16348
rect 9460 16294 9462 16346
rect 9642 16294 9644 16346
rect 9398 16292 9404 16294
rect 9460 16292 9484 16294
rect 9540 16292 9564 16294
rect 9620 16292 9644 16294
rect 9700 16292 9706 16294
rect 9398 16283 9706 16292
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8956 15570 8984 15846
rect 9140 15570 9168 15846
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9398 15260 9706 15269
rect 9398 15258 9404 15260
rect 9460 15258 9484 15260
rect 9540 15258 9564 15260
rect 9620 15258 9644 15260
rect 9700 15258 9706 15260
rect 9460 15206 9462 15258
rect 9642 15206 9644 15258
rect 9398 15204 9404 15206
rect 9460 15204 9484 15206
rect 9540 15204 9564 15206
rect 9620 15204 9644 15206
rect 9700 15204 9706 15206
rect 9398 15195 9706 15204
rect 9398 14172 9706 14181
rect 9398 14170 9404 14172
rect 9460 14170 9484 14172
rect 9540 14170 9564 14172
rect 9620 14170 9644 14172
rect 9700 14170 9706 14172
rect 9460 14118 9462 14170
rect 9642 14118 9644 14170
rect 9398 14116 9404 14118
rect 9460 14116 9484 14118
rect 9540 14116 9564 14118
rect 9620 14116 9644 14118
rect 9700 14116 9706 14118
rect 9398 14107 9706 14116
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12850 8248 13262
rect 9398 13084 9706 13093
rect 9398 13082 9404 13084
rect 9460 13082 9484 13084
rect 9540 13082 9564 13084
rect 9620 13082 9644 13084
rect 9700 13082 9706 13084
rect 9460 13030 9462 13082
rect 9642 13030 9644 13082
rect 9398 13028 9404 13030
rect 9460 13028 9484 13030
rect 9540 13028 9564 13030
rect 9620 13028 9644 13030
rect 9700 13028 9706 13030
rect 9398 13019 9706 13028
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 9398 11996 9706 12005
rect 9398 11994 9404 11996
rect 9460 11994 9484 11996
rect 9540 11994 9564 11996
rect 9620 11994 9644 11996
rect 9700 11994 9706 11996
rect 9460 11942 9462 11994
rect 9642 11942 9644 11994
rect 9398 11940 9404 11942
rect 9460 11940 9484 11942
rect 9540 11940 9564 11942
rect 9620 11940 9644 11942
rect 9700 11940 9706 11942
rect 9398 11931 9706 11940
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9140 10674 9168 11086
rect 9398 10908 9706 10917
rect 9398 10906 9404 10908
rect 9460 10906 9484 10908
rect 9540 10906 9564 10908
rect 9620 10906 9644 10908
rect 9700 10906 9706 10908
rect 9460 10854 9462 10906
rect 9642 10854 9644 10906
rect 9398 10852 9404 10854
rect 9460 10852 9484 10854
rect 9540 10852 9564 10854
rect 9620 10852 9644 10854
rect 9700 10852 9706 10854
rect 9398 10843 9706 10852
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 7852 6886 8156 6914
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4214 7328 4422
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7668 4078 7696 4558
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7852 3942 7880 6886
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7944 4826 7972 5578
rect 8128 5370 8156 6190
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 8220 2854 8248 5034
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5092 1822 5212 1850
rect 5184 800 5212 1822
rect 6472 800 6500 2790
rect 8404 800 8432 5578
rect 8956 2922 8984 10474
rect 9784 10266 9812 10542
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9398 9820 9706 9829
rect 9398 9818 9404 9820
rect 9460 9818 9484 9820
rect 9540 9818 9564 9820
rect 9620 9818 9644 9820
rect 9700 9818 9706 9820
rect 9460 9766 9462 9818
rect 9642 9766 9644 9818
rect 9398 9764 9404 9766
rect 9460 9764 9484 9766
rect 9540 9764 9564 9766
rect 9620 9764 9644 9766
rect 9700 9764 9706 9766
rect 9398 9755 9706 9764
rect 9398 8732 9706 8741
rect 9398 8730 9404 8732
rect 9460 8730 9484 8732
rect 9540 8730 9564 8732
rect 9620 8730 9644 8732
rect 9700 8730 9706 8732
rect 9460 8678 9462 8730
rect 9642 8678 9644 8730
rect 9398 8676 9404 8678
rect 9460 8676 9484 8678
rect 9540 8676 9564 8678
rect 9620 8676 9644 8678
rect 9700 8676 9706 8678
rect 9398 8667 9706 8676
rect 9876 8294 9904 15506
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 13326 10272 15098
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9398 7644 9706 7653
rect 9398 7642 9404 7644
rect 9460 7642 9484 7644
rect 9540 7642 9564 7644
rect 9620 7642 9644 7644
rect 9700 7642 9706 7644
rect 9460 7590 9462 7642
rect 9642 7590 9644 7642
rect 9398 7588 9404 7590
rect 9460 7588 9484 7590
rect 9540 7588 9564 7590
rect 9620 7588 9644 7590
rect 9700 7588 9706 7590
rect 9398 7579 9706 7588
rect 9968 6914 9996 13262
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9784 6886 9996 6914
rect 9784 6798 9812 6886
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9398 6556 9706 6565
rect 9398 6554 9404 6556
rect 9460 6554 9484 6556
rect 9540 6554 9564 6556
rect 9620 6554 9644 6556
rect 9700 6554 9706 6556
rect 9460 6502 9462 6554
rect 9642 6502 9644 6554
rect 9398 6500 9404 6502
rect 9460 6500 9484 6502
rect 9540 6500 9564 6502
rect 9620 6500 9644 6502
rect 9700 6500 9706 6502
rect 9398 6491 9706 6500
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5234 9076 5646
rect 9398 5468 9706 5477
rect 9398 5466 9404 5468
rect 9460 5466 9484 5468
rect 9540 5466 9564 5468
rect 9620 5466 9644 5468
rect 9700 5466 9706 5468
rect 9460 5414 9462 5466
rect 9642 5414 9644 5466
rect 9398 5412 9404 5414
rect 9460 5412 9484 5414
rect 9540 5412 9564 5414
rect 9620 5412 9644 5414
rect 9700 5412 9706 5414
rect 9398 5403 9706 5412
rect 9784 5302 9812 6598
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9398 4380 9706 4389
rect 9398 4378 9404 4380
rect 9460 4378 9484 4380
rect 9540 4378 9564 4380
rect 9620 4378 9644 4380
rect 9700 4378 9706 4380
rect 9460 4326 9462 4378
rect 9642 4326 9644 4378
rect 9398 4324 9404 4326
rect 9460 4324 9484 4326
rect 9540 4324 9564 4326
rect 9620 4324 9644 4326
rect 9700 4324 9706 4326
rect 9398 4315 9706 4324
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3602 9996 3878
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9398 3292 9706 3301
rect 9398 3290 9404 3292
rect 9460 3290 9484 3292
rect 9540 3290 9564 3292
rect 9620 3290 9644 3292
rect 9700 3290 9706 3292
rect 9460 3238 9462 3290
rect 9642 3238 9644 3290
rect 9398 3236 9404 3238
rect 9460 3236 9484 3238
rect 9540 3236 9564 3238
rect 9620 3236 9644 3238
rect 9700 3236 9706 3238
rect 9398 3227 9706 3236
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 9398 2204 9706 2213
rect 9398 2202 9404 2204
rect 9460 2202 9484 2204
rect 9540 2202 9564 2204
rect 9620 2202 9644 2204
rect 9700 2202 9706 2204
rect 9460 2150 9462 2202
rect 9642 2150 9644 2202
rect 9398 2148 9404 2150
rect 9460 2148 9484 2150
rect 9540 2148 9564 2150
rect 9620 2148 9644 2150
rect 9700 2148 9706 2150
rect 9398 2139 9706 2148
rect 9692 870 9904 898
rect 9692 800 9720 870
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 8362 0 8474 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 9876 762 9904 870
rect 10060 762 10088 7754
rect 10336 6914 10364 19314
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18630 10732 18770
rect 11072 18630 11100 24142
rect 13622 23420 13930 23429
rect 13622 23418 13628 23420
rect 13684 23418 13708 23420
rect 13764 23418 13788 23420
rect 13844 23418 13868 23420
rect 13924 23418 13930 23420
rect 13684 23366 13686 23418
rect 13866 23366 13868 23418
rect 13622 23364 13628 23366
rect 13684 23364 13708 23366
rect 13764 23364 13788 23366
rect 13844 23364 13868 23366
rect 13924 23364 13930 23366
rect 13622 23355 13930 23364
rect 13622 22332 13930 22341
rect 13622 22330 13628 22332
rect 13684 22330 13708 22332
rect 13764 22330 13788 22332
rect 13844 22330 13868 22332
rect 13924 22330 13930 22332
rect 13684 22278 13686 22330
rect 13866 22278 13868 22330
rect 13622 22276 13628 22278
rect 13684 22276 13708 22278
rect 13764 22276 13788 22278
rect 13844 22276 13868 22278
rect 13924 22276 13930 22278
rect 13622 22267 13930 22276
rect 13622 21244 13930 21253
rect 13622 21242 13628 21244
rect 13684 21242 13708 21244
rect 13764 21242 13788 21244
rect 13844 21242 13868 21244
rect 13924 21242 13930 21244
rect 13684 21190 13686 21242
rect 13866 21190 13868 21242
rect 13622 21188 13628 21190
rect 13684 21188 13708 21190
rect 13764 21188 13788 21190
rect 13844 21188 13868 21190
rect 13924 21188 13930 21190
rect 13622 21179 13930 21188
rect 13622 20156 13930 20165
rect 13622 20154 13628 20156
rect 13684 20154 13708 20156
rect 13764 20154 13788 20156
rect 13844 20154 13868 20156
rect 13924 20154 13930 20156
rect 13684 20102 13686 20154
rect 13866 20102 13868 20154
rect 13622 20100 13628 20102
rect 13684 20100 13708 20102
rect 13764 20100 13788 20102
rect 13844 20100 13868 20102
rect 13924 20100 13930 20102
rect 13622 20091 13930 20100
rect 16316 20058 16344 29582
rect 17512 26234 17540 36110
rect 17684 36032 17736 36038
rect 17684 35974 17736 35980
rect 17696 35766 17724 35974
rect 17846 35932 18154 35941
rect 17846 35930 17852 35932
rect 17908 35930 17932 35932
rect 17988 35930 18012 35932
rect 18068 35930 18092 35932
rect 18148 35930 18154 35932
rect 17908 35878 17910 35930
rect 18090 35878 18092 35930
rect 17846 35876 17852 35878
rect 17908 35876 17932 35878
rect 17988 35876 18012 35878
rect 18068 35876 18092 35878
rect 18148 35876 18154 35878
rect 17846 35867 18154 35876
rect 17684 35760 17736 35766
rect 17684 35702 17736 35708
rect 19260 35630 19288 39238
rect 19340 38888 19392 38894
rect 19340 38830 19392 38836
rect 19352 38486 19380 38830
rect 19996 38486 20024 41200
rect 19340 38480 19392 38486
rect 19340 38422 19392 38428
rect 19984 38480 20036 38486
rect 19984 38422 20036 38428
rect 20180 38298 20208 41262
rect 20456 41154 20484 41262
rect 20598 41200 20710 42000
rect 21242 41200 21354 42000
rect 21886 41200 21998 42000
rect 22530 41200 22642 42000
rect 23818 41200 23930 42000
rect 24462 41200 24574 42000
rect 25106 41200 25218 42000
rect 25424 41262 25636 41290
rect 20640 41154 20668 41200
rect 20456 41126 20668 41154
rect 22070 39740 22378 39749
rect 22070 39738 22076 39740
rect 22132 39738 22156 39740
rect 22212 39738 22236 39740
rect 22292 39738 22316 39740
rect 22372 39738 22378 39740
rect 22132 39686 22134 39738
rect 22314 39686 22316 39738
rect 22070 39684 22076 39686
rect 22132 39684 22156 39686
rect 22212 39684 22236 39686
rect 22292 39684 22316 39686
rect 22372 39684 22378 39686
rect 22070 39675 22378 39684
rect 20996 39432 21048 39438
rect 20996 39374 21048 39380
rect 22376 39432 22428 39438
rect 22376 39374 22428 39380
rect 20812 39296 20864 39302
rect 20812 39238 20864 39244
rect 20260 38820 20312 38826
rect 20260 38762 20312 38768
rect 19536 38270 20208 38298
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 17846 34844 18154 34853
rect 17846 34842 17852 34844
rect 17908 34842 17932 34844
rect 17988 34842 18012 34844
rect 18068 34842 18092 34844
rect 18148 34842 18154 34844
rect 17908 34790 17910 34842
rect 18090 34790 18092 34842
rect 17846 34788 17852 34790
rect 17908 34788 17932 34790
rect 17988 34788 18012 34790
rect 18068 34788 18092 34790
rect 18148 34788 18154 34790
rect 17846 34779 18154 34788
rect 17846 33756 18154 33765
rect 17846 33754 17852 33756
rect 17908 33754 17932 33756
rect 17988 33754 18012 33756
rect 18068 33754 18092 33756
rect 18148 33754 18154 33756
rect 17908 33702 17910 33754
rect 18090 33702 18092 33754
rect 17846 33700 17852 33702
rect 17908 33700 17932 33702
rect 17988 33700 18012 33702
rect 18068 33700 18092 33702
rect 18148 33700 18154 33702
rect 17846 33691 18154 33700
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 17846 32668 18154 32677
rect 17846 32666 17852 32668
rect 17908 32666 17932 32668
rect 17988 32666 18012 32668
rect 18068 32666 18092 32668
rect 18148 32666 18154 32668
rect 17908 32614 17910 32666
rect 18090 32614 18092 32666
rect 17846 32612 17852 32614
rect 17908 32612 17932 32614
rect 17988 32612 18012 32614
rect 18068 32612 18092 32614
rect 18148 32612 18154 32614
rect 17846 32603 18154 32612
rect 18248 32434 18276 32846
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 17972 32026 18000 32302
rect 17960 32020 18012 32026
rect 17960 31962 18012 31968
rect 19536 31890 19564 38270
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 20088 32502 20116 37878
rect 20272 36854 20300 38762
rect 20824 38282 20852 39238
rect 20904 38888 20956 38894
rect 20904 38830 20956 38836
rect 20812 38276 20864 38282
rect 20812 38218 20864 38224
rect 20916 38010 20944 38830
rect 21008 38418 21036 39374
rect 21088 39364 21140 39370
rect 21088 39306 21140 39312
rect 21100 38962 21128 39306
rect 22388 38962 22416 39374
rect 22572 39250 22600 41200
rect 22572 39222 22692 39250
rect 21088 38956 21140 38962
rect 21088 38898 21140 38904
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22070 38652 22378 38661
rect 22070 38650 22076 38652
rect 22132 38650 22156 38652
rect 22212 38650 22236 38652
rect 22292 38650 22316 38652
rect 22372 38650 22378 38652
rect 22132 38598 22134 38650
rect 22314 38598 22316 38650
rect 22070 38596 22076 38598
rect 22132 38596 22156 38598
rect 22212 38596 22236 38598
rect 22292 38596 22316 38598
rect 22372 38596 22378 38598
rect 22070 38587 22378 38596
rect 22572 38554 22600 38830
rect 22560 38548 22612 38554
rect 22560 38490 22612 38496
rect 20996 38412 21048 38418
rect 20996 38354 21048 38360
rect 20904 38004 20956 38010
rect 20904 37946 20956 37952
rect 22468 37664 22520 37670
rect 22468 37606 22520 37612
rect 22070 37564 22378 37573
rect 22070 37562 22076 37564
rect 22132 37562 22156 37564
rect 22212 37562 22236 37564
rect 22292 37562 22316 37564
rect 22372 37562 22378 37564
rect 22132 37510 22134 37562
rect 22314 37510 22316 37562
rect 22070 37508 22076 37510
rect 22132 37508 22156 37510
rect 22212 37508 22236 37510
rect 22292 37508 22316 37510
rect 22372 37508 22378 37510
rect 22070 37499 22378 37508
rect 22480 37330 22508 37606
rect 22664 37330 22692 39222
rect 25148 39030 25176 41200
rect 25136 39024 25188 39030
rect 25136 38966 25188 38972
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 22468 37324 22520 37330
rect 22468 37266 22520 37272
rect 22652 37324 22704 37330
rect 22652 37266 22704 37272
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 22204 36922 22232 37130
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 20260 36848 20312 36854
rect 20260 36790 20312 36796
rect 22070 36476 22378 36485
rect 22070 36474 22076 36476
rect 22132 36474 22156 36476
rect 22212 36474 22236 36476
rect 22292 36474 22316 36476
rect 22372 36474 22378 36476
rect 22132 36422 22134 36474
rect 22314 36422 22316 36474
rect 22070 36420 22076 36422
rect 22132 36420 22156 36422
rect 22212 36420 22236 36422
rect 22292 36420 22316 36422
rect 22372 36420 22378 36422
rect 22070 36411 22378 36420
rect 22070 35388 22378 35397
rect 22070 35386 22076 35388
rect 22132 35386 22156 35388
rect 22212 35386 22236 35388
rect 22292 35386 22316 35388
rect 22372 35386 22378 35388
rect 22132 35334 22134 35386
rect 22314 35334 22316 35386
rect 22070 35332 22076 35334
rect 22132 35332 22156 35334
rect 22212 35332 22236 35334
rect 22292 35332 22316 35334
rect 22372 35332 22378 35334
rect 22070 35323 22378 35332
rect 22070 34300 22378 34309
rect 22070 34298 22076 34300
rect 22132 34298 22156 34300
rect 22212 34298 22236 34300
rect 22292 34298 22316 34300
rect 22372 34298 22378 34300
rect 22132 34246 22134 34298
rect 22314 34246 22316 34298
rect 22070 34244 22076 34246
rect 22132 34244 22156 34246
rect 22212 34244 22236 34246
rect 22292 34244 22316 34246
rect 22372 34244 22378 34246
rect 22070 34235 22378 34244
rect 22070 33212 22378 33221
rect 22070 33210 22076 33212
rect 22132 33210 22156 33212
rect 22212 33210 22236 33212
rect 22292 33210 22316 33212
rect 22372 33210 22378 33212
rect 22132 33158 22134 33210
rect 22314 33158 22316 33210
rect 22070 33156 22076 33158
rect 22132 33156 22156 33158
rect 22212 33156 22236 33158
rect 22292 33156 22316 33158
rect 22372 33156 22378 33158
rect 22070 33147 22378 33156
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 22070 32124 22378 32133
rect 22070 32122 22076 32124
rect 22132 32122 22156 32124
rect 22212 32122 22236 32124
rect 22292 32122 22316 32124
rect 22372 32122 22378 32124
rect 22132 32070 22134 32122
rect 22314 32070 22316 32122
rect 22070 32068 22076 32070
rect 22132 32068 22156 32070
rect 22212 32068 22236 32070
rect 22292 32068 22316 32070
rect 22372 32068 22378 32070
rect 22070 32059 22378 32068
rect 17592 31884 17644 31890
rect 17592 31826 17644 31832
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 17328 26206 17540 26234
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16592 20466 16620 23666
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 19514 11652 19722
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 13622 19068 13930 19077
rect 13622 19066 13628 19068
rect 13684 19066 13708 19068
rect 13764 19066 13788 19068
rect 13844 19066 13868 19068
rect 13924 19066 13930 19068
rect 13684 19014 13686 19066
rect 13866 19014 13868 19066
rect 13622 19012 13628 19014
rect 13684 19012 13708 19014
rect 13764 19012 13788 19014
rect 13844 19012 13868 19014
rect 13924 19012 13930 19014
rect 13622 19003 13930 19012
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 13622 17980 13930 17989
rect 13622 17978 13628 17980
rect 13684 17978 13708 17980
rect 13764 17978 13788 17980
rect 13844 17978 13868 17980
rect 13924 17978 13930 17980
rect 13684 17926 13686 17978
rect 13866 17926 13868 17978
rect 13622 17924 13628 17926
rect 13684 17924 13708 17926
rect 13764 17924 13788 17926
rect 13844 17924 13868 17926
rect 13924 17924 13930 17926
rect 13622 17915 13930 17924
rect 13622 16892 13930 16901
rect 13622 16890 13628 16892
rect 13684 16890 13708 16892
rect 13764 16890 13788 16892
rect 13844 16890 13868 16892
rect 13924 16890 13930 16892
rect 13684 16838 13686 16890
rect 13866 16838 13868 16890
rect 13622 16836 13628 16838
rect 13684 16836 13708 16838
rect 13764 16836 13788 16838
rect 13844 16836 13868 16838
rect 13924 16836 13930 16838
rect 13622 16827 13930 16836
rect 13622 15804 13930 15813
rect 13622 15802 13628 15804
rect 13684 15802 13708 15804
rect 13764 15802 13788 15804
rect 13844 15802 13868 15804
rect 13924 15802 13930 15804
rect 13684 15750 13686 15802
rect 13866 15750 13868 15802
rect 13622 15748 13628 15750
rect 13684 15748 13708 15750
rect 13764 15748 13788 15750
rect 13844 15748 13868 15750
rect 13924 15748 13930 15750
rect 13622 15739 13930 15748
rect 13622 14716 13930 14725
rect 13622 14714 13628 14716
rect 13684 14714 13708 14716
rect 13764 14714 13788 14716
rect 13844 14714 13868 14716
rect 13924 14714 13930 14716
rect 13684 14662 13686 14714
rect 13866 14662 13868 14714
rect 13622 14660 13628 14662
rect 13684 14660 13708 14662
rect 13764 14660 13788 14662
rect 13844 14660 13868 14662
rect 13924 14660 13930 14662
rect 13622 14651 13930 14660
rect 13622 13628 13930 13637
rect 13622 13626 13628 13628
rect 13684 13626 13708 13628
rect 13764 13626 13788 13628
rect 13844 13626 13868 13628
rect 13924 13626 13930 13628
rect 13684 13574 13686 13626
rect 13866 13574 13868 13626
rect 13622 13572 13628 13574
rect 13684 13572 13708 13574
rect 13764 13572 13788 13574
rect 13844 13572 13868 13574
rect 13924 13572 13930 13574
rect 13622 13563 13930 13572
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 10130 10456 13126
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14384 12646 14412 12922
rect 16316 12646 16344 19994
rect 16868 19786 16896 20198
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16868 19378 16896 19722
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 13622 12540 13930 12549
rect 13622 12538 13628 12540
rect 13684 12538 13708 12540
rect 13764 12538 13788 12540
rect 13844 12538 13868 12540
rect 13924 12538 13930 12540
rect 13684 12486 13686 12538
rect 13866 12486 13868 12538
rect 13622 12484 13628 12486
rect 13684 12484 13708 12486
rect 13764 12484 13788 12486
rect 13844 12484 13868 12486
rect 13924 12484 13930 12486
rect 13622 12475 13930 12484
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 13622 11452 13930 11461
rect 13622 11450 13628 11452
rect 13684 11450 13708 11452
rect 13764 11450 13788 11452
rect 13844 11450 13868 11452
rect 13924 11450 13930 11452
rect 13684 11398 13686 11450
rect 13866 11398 13868 11450
rect 13622 11396 13628 11398
rect 13684 11396 13708 11398
rect 13764 11396 13788 11398
rect 13844 11396 13868 11398
rect 13924 11396 13930 11398
rect 13622 11387 13930 11396
rect 14292 11218 14320 11494
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14384 10674 14412 12582
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14476 10810 14504 11018
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 13622 10364 13930 10373
rect 13622 10362 13628 10364
rect 13684 10362 13708 10364
rect 13764 10362 13788 10364
rect 13844 10362 13868 10364
rect 13924 10362 13930 10364
rect 13684 10310 13686 10362
rect 13866 10310 13868 10362
rect 13622 10308 13628 10310
rect 13684 10308 13708 10310
rect 13764 10308 13788 10310
rect 13844 10308 13868 10310
rect 13924 10308 13930 10310
rect 13622 10299 13930 10308
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 9586 11928 9998
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9654 12112 9862
rect 12176 9654 12204 9930
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 12176 8498 12204 9590
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 7954 12940 8366
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13096 7954 13124 8298
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 10244 6886 10364 6914
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 5778 10180 6734
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10244 3738 10272 6886
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 6322 12848 6734
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6390 13032 6598
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5778 10364 6054
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5370 10640 5714
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10704 5166 10732 6258
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11164 4690 11192 4966
rect 11624 4758 11652 4966
rect 13280 4826 13308 6190
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10520 3670 10548 3878
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10336 800 10364 3538
rect 13464 2582 13492 9454
rect 13622 9276 13930 9285
rect 13622 9274 13628 9276
rect 13684 9274 13708 9276
rect 13764 9274 13788 9276
rect 13844 9274 13868 9276
rect 13924 9274 13930 9276
rect 13684 9222 13686 9274
rect 13866 9222 13868 9274
rect 13622 9220 13628 9222
rect 13684 9220 13708 9222
rect 13764 9220 13788 9222
rect 13844 9220 13868 9222
rect 13924 9220 13930 9222
rect 13622 9211 13930 9220
rect 13622 8188 13930 8197
rect 13622 8186 13628 8188
rect 13684 8186 13708 8188
rect 13764 8186 13788 8188
rect 13844 8186 13868 8188
rect 13924 8186 13930 8188
rect 13684 8134 13686 8186
rect 13866 8134 13868 8186
rect 13622 8132 13628 8134
rect 13684 8132 13708 8134
rect 13764 8132 13788 8134
rect 13844 8132 13868 8134
rect 13924 8132 13930 8134
rect 13622 8123 13930 8132
rect 13622 7100 13930 7109
rect 13622 7098 13628 7100
rect 13684 7098 13708 7100
rect 13764 7098 13788 7100
rect 13844 7098 13868 7100
rect 13924 7098 13930 7100
rect 13684 7046 13686 7098
rect 13866 7046 13868 7098
rect 13622 7044 13628 7046
rect 13684 7044 13708 7046
rect 13764 7044 13788 7046
rect 13844 7044 13868 7046
rect 13924 7044 13930 7046
rect 13622 7035 13930 7044
rect 13622 6012 13930 6021
rect 13622 6010 13628 6012
rect 13684 6010 13708 6012
rect 13764 6010 13788 6012
rect 13844 6010 13868 6012
rect 13924 6010 13930 6012
rect 13684 5958 13686 6010
rect 13866 5958 13868 6010
rect 13622 5956 13628 5958
rect 13684 5956 13708 5958
rect 13764 5956 13788 5958
rect 13844 5956 13868 5958
rect 13924 5956 13930 5958
rect 13622 5947 13930 5956
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13556 800 13584 5578
rect 13622 4924 13930 4933
rect 13622 4922 13628 4924
rect 13684 4922 13708 4924
rect 13764 4922 13788 4924
rect 13844 4922 13868 4924
rect 13924 4922 13930 4924
rect 13684 4870 13686 4922
rect 13866 4870 13868 4922
rect 13622 4868 13628 4870
rect 13684 4868 13708 4870
rect 13764 4868 13788 4870
rect 13844 4868 13868 4870
rect 13924 4868 13930 4870
rect 13622 4859 13930 4868
rect 13622 3836 13930 3845
rect 13622 3834 13628 3836
rect 13684 3834 13708 3836
rect 13764 3834 13788 3836
rect 13844 3834 13868 3836
rect 13924 3834 13930 3836
rect 13684 3782 13686 3834
rect 13866 3782 13868 3834
rect 13622 3780 13628 3782
rect 13684 3780 13708 3782
rect 13764 3780 13788 3782
rect 13844 3780 13868 3782
rect 13924 3780 13930 3782
rect 13622 3771 13930 3780
rect 13622 2748 13930 2757
rect 13622 2746 13628 2748
rect 13684 2746 13708 2748
rect 13764 2746 13788 2748
rect 13844 2746 13868 2748
rect 13924 2746 13930 2748
rect 13684 2694 13686 2746
rect 13866 2694 13868 2746
rect 13622 2692 13628 2694
rect 13684 2692 13708 2694
rect 13764 2692 13788 2694
rect 13844 2692 13868 2694
rect 13924 2692 13930 2694
rect 13622 2683 13930 2692
rect 14844 800 14872 11154
rect 16500 10062 16528 18566
rect 16960 18426 16988 21422
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20466 17264 20878
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17052 19922 17080 20402
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17052 16574 17080 19246
rect 17144 18086 17172 19382
rect 17236 18766 17264 20402
rect 17328 18970 17356 26206
rect 17604 20806 17632 31826
rect 20260 31748 20312 31754
rect 20260 31690 20312 31696
rect 17846 31580 18154 31589
rect 17846 31578 17852 31580
rect 17908 31578 17932 31580
rect 17988 31578 18012 31580
rect 18068 31578 18092 31580
rect 18148 31578 18154 31580
rect 17908 31526 17910 31578
rect 18090 31526 18092 31578
rect 17846 31524 17852 31526
rect 17908 31524 17932 31526
rect 17988 31524 18012 31526
rect 18068 31524 18092 31526
rect 18148 31524 18154 31526
rect 17846 31515 18154 31524
rect 20272 31482 20300 31690
rect 20260 31476 20312 31482
rect 20260 31418 20312 31424
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 17846 30492 18154 30501
rect 17846 30490 17852 30492
rect 17908 30490 17932 30492
rect 17988 30490 18012 30492
rect 18068 30490 18092 30492
rect 18148 30490 18154 30492
rect 17908 30438 17910 30490
rect 18090 30438 18092 30490
rect 17846 30436 17852 30438
rect 17908 30436 17932 30438
rect 17988 30436 18012 30438
rect 18068 30436 18092 30438
rect 18148 30436 18154 30438
rect 17846 30427 18154 30436
rect 17846 29404 18154 29413
rect 17846 29402 17852 29404
rect 17908 29402 17932 29404
rect 17988 29402 18012 29404
rect 18068 29402 18092 29404
rect 18148 29402 18154 29404
rect 17908 29350 17910 29402
rect 18090 29350 18092 29402
rect 17846 29348 17852 29350
rect 17908 29348 17932 29350
rect 17988 29348 18012 29350
rect 18068 29348 18092 29350
rect 18148 29348 18154 29350
rect 17846 29339 18154 29348
rect 17846 28316 18154 28325
rect 17846 28314 17852 28316
rect 17908 28314 17932 28316
rect 17988 28314 18012 28316
rect 18068 28314 18092 28316
rect 18148 28314 18154 28316
rect 17908 28262 17910 28314
rect 18090 28262 18092 28314
rect 17846 28260 17852 28262
rect 17908 28260 17932 28262
rect 17988 28260 18012 28262
rect 18068 28260 18092 28262
rect 18148 28260 18154 28262
rect 17846 28251 18154 28260
rect 17846 27228 18154 27237
rect 17846 27226 17852 27228
rect 17908 27226 17932 27228
rect 17988 27226 18012 27228
rect 18068 27226 18092 27228
rect 18148 27226 18154 27228
rect 17908 27174 17910 27226
rect 18090 27174 18092 27226
rect 17846 27172 17852 27174
rect 17908 27172 17932 27174
rect 17988 27172 18012 27174
rect 18068 27172 18092 27174
rect 18148 27172 18154 27174
rect 17846 27163 18154 27172
rect 17846 26140 18154 26149
rect 17846 26138 17852 26140
rect 17908 26138 17932 26140
rect 17988 26138 18012 26140
rect 18068 26138 18092 26140
rect 18148 26138 18154 26140
rect 17908 26086 17910 26138
rect 18090 26086 18092 26138
rect 17846 26084 17852 26086
rect 17908 26084 17932 26086
rect 17988 26084 18012 26086
rect 18068 26084 18092 26086
rect 18148 26084 18154 26086
rect 17846 26075 18154 26084
rect 17846 25052 18154 25061
rect 17846 25050 17852 25052
rect 17908 25050 17932 25052
rect 17988 25050 18012 25052
rect 18068 25050 18092 25052
rect 18148 25050 18154 25052
rect 17908 24998 17910 25050
rect 18090 24998 18092 25050
rect 17846 24996 17852 24998
rect 17908 24996 17932 24998
rect 17988 24996 18012 24998
rect 18068 24996 18092 24998
rect 18148 24996 18154 24998
rect 17846 24987 18154 24996
rect 17846 23964 18154 23973
rect 17846 23962 17852 23964
rect 17908 23962 17932 23964
rect 17988 23962 18012 23964
rect 18068 23962 18092 23964
rect 18148 23962 18154 23964
rect 17908 23910 17910 23962
rect 18090 23910 18092 23962
rect 17846 23908 17852 23910
rect 17908 23908 17932 23910
rect 17988 23908 18012 23910
rect 18068 23908 18092 23910
rect 18148 23908 18154 23910
rect 17846 23899 18154 23908
rect 17846 22876 18154 22885
rect 17846 22874 17852 22876
rect 17908 22874 17932 22876
rect 17988 22874 18012 22876
rect 18068 22874 18092 22876
rect 18148 22874 18154 22876
rect 17908 22822 17910 22874
rect 18090 22822 18092 22874
rect 17846 22820 17852 22822
rect 17908 22820 17932 22822
rect 17988 22820 18012 22822
rect 18068 22820 18092 22822
rect 18148 22820 18154 22822
rect 17846 22811 18154 22820
rect 17846 21788 18154 21797
rect 17846 21786 17852 21788
rect 17908 21786 17932 21788
rect 17988 21786 18012 21788
rect 18068 21786 18092 21788
rect 18148 21786 18154 21788
rect 17908 21734 17910 21786
rect 18090 21734 18092 21786
rect 17846 21732 17852 21734
rect 17908 21732 17932 21734
rect 17988 21732 18012 21734
rect 18068 21732 18092 21734
rect 18148 21732 18154 21734
rect 17846 21723 18154 21732
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17696 20942 17724 21490
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 19990 17632 20742
rect 17846 20700 18154 20709
rect 17846 20698 17852 20700
rect 17908 20698 17932 20700
rect 17988 20698 18012 20700
rect 18068 20698 18092 20700
rect 18148 20698 18154 20700
rect 17908 20646 17910 20698
rect 18090 20646 18092 20698
rect 17846 20644 17852 20646
rect 17908 20644 17932 20646
rect 17988 20644 18012 20646
rect 18068 20644 18092 20646
rect 18148 20644 18154 20646
rect 17846 20635 18154 20644
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19378 17448 19790
rect 17846 19612 18154 19621
rect 17846 19610 17852 19612
rect 17908 19610 17932 19612
rect 17988 19610 18012 19612
rect 18068 19610 18092 19612
rect 18148 19610 18154 19612
rect 17908 19558 17910 19610
rect 18090 19558 18092 19610
rect 17846 19556 17852 19558
rect 17908 19556 17932 19558
rect 17988 19556 18012 19558
rect 18068 19556 18092 19558
rect 18148 19556 18154 19558
rect 17846 19547 18154 19556
rect 18248 19446 18276 30602
rect 20180 30394 20208 31282
rect 22070 31036 22378 31045
rect 22070 31034 22076 31036
rect 22132 31034 22156 31036
rect 22212 31034 22236 31036
rect 22292 31034 22316 31036
rect 22372 31034 22378 31036
rect 22132 30982 22134 31034
rect 22314 30982 22316 31034
rect 22070 30980 22076 30982
rect 22132 30980 22156 30982
rect 22212 30980 22236 30982
rect 22292 30980 22316 30982
rect 22372 30980 22378 30982
rect 22070 30971 22378 30980
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19352 29714 19380 29990
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 18340 24818 18368 29242
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 23798 18368 24754
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 19352 23526 19380 29446
rect 19812 29306 19840 29514
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19708 28552 19760 28558
rect 19708 28494 19760 28500
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19628 23730 19656 24074
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17236 18358 17264 18702
rect 17420 18698 17448 19314
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16684 16546 17080 16574
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16684 9926 16712 16546
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16500 9654 16528 9862
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16776 6914 16804 13398
rect 16868 13394 16896 13670
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11218 16896 11494
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16776 6886 16896 6914
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 5778 15792 6598
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5778 15976 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3058 15608 3470
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15764 2650 15792 3402
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16132 800 16160 3538
rect 16868 2258 16896 6886
rect 16960 3058 16988 15846
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13394 17080 13670
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11218 17080 11494
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17144 6390 17172 18022
rect 17420 16182 17448 18634
rect 17512 18290 17540 19178
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17604 17678 17632 18294
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17420 15502 17448 16118
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17512 15162 17540 15302
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17696 13938 17724 18906
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17696 10742 17724 13874
rect 17788 11762 17816 18566
rect 17846 18524 18154 18533
rect 17846 18522 17852 18524
rect 17908 18522 17932 18524
rect 17988 18522 18012 18524
rect 18068 18522 18092 18524
rect 18148 18522 18154 18524
rect 17908 18470 17910 18522
rect 18090 18470 18092 18522
rect 17846 18468 17852 18470
rect 17908 18468 17932 18470
rect 17988 18468 18012 18470
rect 18068 18468 18092 18470
rect 18148 18468 18154 18470
rect 17846 18459 18154 18468
rect 17846 17436 18154 17445
rect 17846 17434 17852 17436
rect 17908 17434 17932 17436
rect 17988 17434 18012 17436
rect 18068 17434 18092 17436
rect 18148 17434 18154 17436
rect 17908 17382 17910 17434
rect 18090 17382 18092 17434
rect 17846 17380 17852 17382
rect 17908 17380 17932 17382
rect 17988 17380 18012 17382
rect 18068 17380 18092 17382
rect 18148 17380 18154 17382
rect 17846 17371 18154 17380
rect 17846 16348 18154 16357
rect 17846 16346 17852 16348
rect 17908 16346 17932 16348
rect 17988 16346 18012 16348
rect 18068 16346 18092 16348
rect 18148 16346 18154 16348
rect 17908 16294 17910 16346
rect 18090 16294 18092 16346
rect 17846 16292 17852 16294
rect 17908 16292 17932 16294
rect 17988 16292 18012 16294
rect 18068 16292 18092 16294
rect 18148 16292 18154 16294
rect 17846 16283 18154 16292
rect 18248 16182 18276 19382
rect 18708 19378 18736 20402
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 17846 15260 18154 15269
rect 17846 15258 17852 15260
rect 17908 15258 17932 15260
rect 17988 15258 18012 15260
rect 18068 15258 18092 15260
rect 18148 15258 18154 15260
rect 17908 15206 17910 15258
rect 18090 15206 18092 15258
rect 17846 15204 17852 15206
rect 17908 15204 17932 15206
rect 17988 15204 18012 15206
rect 18068 15204 18092 15206
rect 18148 15204 18154 15206
rect 17846 15195 18154 15204
rect 17846 14172 18154 14181
rect 17846 14170 17852 14172
rect 17908 14170 17932 14172
rect 17988 14170 18012 14172
rect 18068 14170 18092 14172
rect 18148 14170 18154 14172
rect 17908 14118 17910 14170
rect 18090 14118 18092 14170
rect 17846 14116 17852 14118
rect 17908 14116 17932 14118
rect 17988 14116 18012 14118
rect 18068 14116 18092 14118
rect 18148 14116 18154 14118
rect 17846 14107 18154 14116
rect 17846 13084 18154 13093
rect 17846 13082 17852 13084
rect 17908 13082 17932 13084
rect 17988 13082 18012 13084
rect 18068 13082 18092 13084
rect 18148 13082 18154 13084
rect 17908 13030 17910 13082
rect 18090 13030 18092 13082
rect 17846 13028 17852 13030
rect 17908 13028 17932 13030
rect 17988 13028 18012 13030
rect 18068 13028 18092 13030
rect 18148 13028 18154 13030
rect 17846 13019 18154 13028
rect 17846 11996 18154 12005
rect 17846 11994 17852 11996
rect 17908 11994 17932 11996
rect 17988 11994 18012 11996
rect 18068 11994 18092 11996
rect 18148 11994 18154 11996
rect 17908 11942 17910 11994
rect 18090 11942 18092 11994
rect 17846 11940 17852 11942
rect 17908 11940 17932 11942
rect 17988 11940 18012 11942
rect 18068 11940 18092 11942
rect 18148 11940 18154 11942
rect 17846 11931 18154 11940
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17846 10908 18154 10917
rect 17846 10906 17852 10908
rect 17908 10906 17932 10908
rect 17988 10906 18012 10908
rect 18068 10906 18092 10908
rect 18148 10906 18154 10908
rect 17908 10854 17910 10906
rect 18090 10854 18092 10906
rect 17846 10852 17852 10854
rect 17908 10852 17932 10854
rect 17988 10852 18012 10854
rect 18068 10852 18092 10854
rect 18148 10852 18154 10854
rect 17846 10843 18154 10852
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17846 9820 18154 9829
rect 17846 9818 17852 9820
rect 17908 9818 17932 9820
rect 17988 9818 18012 9820
rect 18068 9818 18092 9820
rect 18148 9818 18154 9820
rect 17908 9766 17910 9818
rect 18090 9766 18092 9818
rect 17846 9764 17852 9766
rect 17908 9764 17932 9766
rect 17988 9764 18012 9766
rect 18068 9764 18092 9766
rect 18148 9764 18154 9766
rect 17846 9755 18154 9764
rect 17846 8732 18154 8741
rect 17846 8730 17852 8732
rect 17908 8730 17932 8732
rect 17988 8730 18012 8732
rect 18068 8730 18092 8732
rect 18148 8730 18154 8732
rect 17908 8678 17910 8730
rect 18090 8678 18092 8730
rect 17846 8676 17852 8678
rect 17908 8676 17932 8678
rect 17988 8676 18012 8678
rect 18068 8676 18092 8678
rect 18148 8676 18154 8678
rect 17846 8667 18154 8676
rect 17846 7644 18154 7653
rect 17846 7642 17852 7644
rect 17908 7642 17932 7644
rect 17988 7642 18012 7644
rect 18068 7642 18092 7644
rect 18148 7642 18154 7644
rect 17908 7590 17910 7642
rect 18090 7590 18092 7642
rect 17846 7588 17852 7590
rect 17908 7588 17932 7590
rect 17988 7588 18012 7590
rect 18068 7588 18092 7590
rect 18148 7588 18154 7590
rect 17846 7579 18154 7588
rect 17846 6556 18154 6565
rect 17846 6554 17852 6556
rect 17908 6554 17932 6556
rect 17988 6554 18012 6556
rect 18068 6554 18092 6556
rect 18148 6554 18154 6556
rect 17908 6502 17910 6554
rect 18090 6502 18092 6554
rect 17846 6500 17852 6502
rect 17908 6500 17932 6502
rect 17988 6500 18012 6502
rect 18068 6500 18092 6502
rect 18148 6500 18154 6502
rect 17846 6491 18154 6500
rect 18892 6458 18920 19382
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 15366 19012 15438
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18984 15026 19012 15302
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19168 14958 19196 18838
rect 19352 18834 19380 23462
rect 19720 22982 19748 28494
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19996 23118 20024 23666
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19628 9654 19656 9862
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19444 9178 19472 9454
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19720 6798 19748 22918
rect 20180 19514 20208 30330
rect 22070 29948 22378 29957
rect 22070 29946 22076 29948
rect 22132 29946 22156 29948
rect 22212 29946 22236 29948
rect 22292 29946 22316 29948
rect 22372 29946 22378 29948
rect 22132 29894 22134 29946
rect 22314 29894 22316 29946
rect 22070 29892 22076 29894
rect 22132 29892 22156 29894
rect 22212 29892 22236 29894
rect 22292 29892 22316 29894
rect 22372 29892 22378 29894
rect 22070 29883 22378 29892
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 29170 20760 29446
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20732 23526 20760 29106
rect 22070 28860 22378 28869
rect 22070 28858 22076 28860
rect 22132 28858 22156 28860
rect 22212 28858 22236 28860
rect 22292 28858 22316 28860
rect 22372 28858 22378 28860
rect 22132 28806 22134 28858
rect 22314 28806 22316 28858
rect 22070 28804 22076 28806
rect 22132 28804 22156 28806
rect 22212 28804 22236 28806
rect 22292 28804 22316 28806
rect 22372 28804 22378 28806
rect 22070 28795 22378 28804
rect 22070 27772 22378 27781
rect 22070 27770 22076 27772
rect 22132 27770 22156 27772
rect 22212 27770 22236 27772
rect 22292 27770 22316 27772
rect 22372 27770 22378 27772
rect 22132 27718 22134 27770
rect 22314 27718 22316 27770
rect 22070 27716 22076 27718
rect 22132 27716 22156 27718
rect 22212 27716 22236 27718
rect 22292 27716 22316 27718
rect 22372 27716 22378 27718
rect 22070 27707 22378 27716
rect 22070 26684 22378 26693
rect 22070 26682 22076 26684
rect 22132 26682 22156 26684
rect 22212 26682 22236 26684
rect 22292 26682 22316 26684
rect 22372 26682 22378 26684
rect 22132 26630 22134 26682
rect 22314 26630 22316 26682
rect 22070 26628 22076 26630
rect 22132 26628 22156 26630
rect 22212 26628 22236 26630
rect 22292 26628 22316 26630
rect 22372 26628 22378 26630
rect 22070 26619 22378 26628
rect 22070 25596 22378 25605
rect 22070 25594 22076 25596
rect 22132 25594 22156 25596
rect 22212 25594 22236 25596
rect 22292 25594 22316 25596
rect 22372 25594 22378 25596
rect 22132 25542 22134 25594
rect 22314 25542 22316 25594
rect 22070 25540 22076 25542
rect 22132 25540 22156 25542
rect 22212 25540 22236 25542
rect 22292 25540 22316 25542
rect 22372 25540 22378 25542
rect 22070 25531 22378 25540
rect 22070 24508 22378 24517
rect 22070 24506 22076 24508
rect 22132 24506 22156 24508
rect 22212 24506 22236 24508
rect 22292 24506 22316 24508
rect 22372 24506 22378 24508
rect 22132 24454 22134 24506
rect 22314 24454 22316 24506
rect 22070 24452 22076 24454
rect 22132 24452 22156 24454
rect 22212 24452 22236 24454
rect 22292 24452 22316 24454
rect 22372 24452 22378 24454
rect 22070 24443 22378 24452
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20732 20466 20760 23462
rect 22070 23420 22378 23429
rect 22070 23418 22076 23420
rect 22132 23418 22156 23420
rect 22212 23418 22236 23420
rect 22292 23418 22316 23420
rect 22372 23418 22378 23420
rect 22132 23366 22134 23418
rect 22314 23366 22316 23418
rect 22070 23364 22076 23366
rect 22132 23364 22156 23366
rect 22212 23364 22236 23366
rect 22292 23364 22316 23366
rect 22372 23364 22378 23366
rect 22070 23355 22378 23364
rect 22070 22332 22378 22341
rect 22070 22330 22076 22332
rect 22132 22330 22156 22332
rect 22212 22330 22236 22332
rect 22292 22330 22316 22332
rect 22372 22330 22378 22332
rect 22132 22278 22134 22330
rect 22314 22278 22316 22330
rect 22070 22276 22076 22278
rect 22132 22276 22156 22278
rect 22212 22276 22236 22278
rect 22292 22276 22316 22278
rect 22372 22276 22378 22278
rect 22070 22267 22378 22276
rect 23492 21486 23520 38286
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24872 28558 24900 31282
rect 25424 29714 25452 41262
rect 25608 41154 25636 41262
rect 25750 41200 25862 42000
rect 26394 41200 26506 42000
rect 26712 41262 26924 41290
rect 25792 41154 25820 41200
rect 25608 41126 25820 41154
rect 26294 39196 26602 39205
rect 26294 39194 26300 39196
rect 26356 39194 26380 39196
rect 26436 39194 26460 39196
rect 26516 39194 26540 39196
rect 26596 39194 26602 39196
rect 26356 39142 26358 39194
rect 26538 39142 26540 39194
rect 26294 39140 26300 39142
rect 26356 39140 26380 39142
rect 26436 39140 26460 39142
rect 26516 39140 26540 39142
rect 26596 39140 26602 39142
rect 26294 39131 26602 39140
rect 26294 38108 26602 38117
rect 26294 38106 26300 38108
rect 26356 38106 26380 38108
rect 26436 38106 26460 38108
rect 26516 38106 26540 38108
rect 26596 38106 26602 38108
rect 26356 38054 26358 38106
rect 26538 38054 26540 38106
rect 26294 38052 26300 38054
rect 26356 38052 26380 38054
rect 26436 38052 26460 38054
rect 26516 38052 26540 38054
rect 26596 38052 26602 38054
rect 26294 38043 26602 38052
rect 26294 37020 26602 37029
rect 26294 37018 26300 37020
rect 26356 37018 26380 37020
rect 26436 37018 26460 37020
rect 26516 37018 26540 37020
rect 26596 37018 26602 37020
rect 26356 36966 26358 37018
rect 26538 36966 26540 37018
rect 26294 36964 26300 36966
rect 26356 36964 26380 36966
rect 26436 36964 26460 36966
rect 26516 36964 26540 36966
rect 26596 36964 26602 36966
rect 26294 36955 26602 36964
rect 26294 35932 26602 35941
rect 26294 35930 26300 35932
rect 26356 35930 26380 35932
rect 26436 35930 26460 35932
rect 26516 35930 26540 35932
rect 26596 35930 26602 35932
rect 26356 35878 26358 35930
rect 26538 35878 26540 35930
rect 26294 35876 26300 35878
rect 26356 35876 26380 35878
rect 26436 35876 26460 35878
rect 26516 35876 26540 35878
rect 26596 35876 26602 35878
rect 26294 35867 26602 35876
rect 26294 34844 26602 34853
rect 26294 34842 26300 34844
rect 26356 34842 26380 34844
rect 26436 34842 26460 34844
rect 26516 34842 26540 34844
rect 26596 34842 26602 34844
rect 26356 34790 26358 34842
rect 26538 34790 26540 34842
rect 26294 34788 26300 34790
rect 26356 34788 26380 34790
rect 26436 34788 26460 34790
rect 26516 34788 26540 34790
rect 26596 34788 26602 34790
rect 26294 34779 26602 34788
rect 26294 33756 26602 33765
rect 26294 33754 26300 33756
rect 26356 33754 26380 33756
rect 26436 33754 26460 33756
rect 26516 33754 26540 33756
rect 26596 33754 26602 33756
rect 26356 33702 26358 33754
rect 26538 33702 26540 33754
rect 26294 33700 26300 33702
rect 26356 33700 26380 33702
rect 26436 33700 26460 33702
rect 26516 33700 26540 33702
rect 26596 33700 26602 33702
rect 26294 33691 26602 33700
rect 26294 32668 26602 32677
rect 26294 32666 26300 32668
rect 26356 32666 26380 32668
rect 26436 32666 26460 32668
rect 26516 32666 26540 32668
rect 26596 32666 26602 32668
rect 26356 32614 26358 32666
rect 26538 32614 26540 32666
rect 26294 32612 26300 32614
rect 26356 32612 26380 32614
rect 26436 32612 26460 32614
rect 26516 32612 26540 32614
rect 26596 32612 26602 32614
rect 26294 32603 26602 32612
rect 26294 31580 26602 31589
rect 26294 31578 26300 31580
rect 26356 31578 26380 31580
rect 26436 31578 26460 31580
rect 26516 31578 26540 31580
rect 26596 31578 26602 31580
rect 26356 31526 26358 31578
rect 26538 31526 26540 31578
rect 26294 31524 26300 31526
rect 26356 31524 26380 31526
rect 26436 31524 26460 31526
rect 26516 31524 26540 31526
rect 26596 31524 26602 31526
rect 26294 31515 26602 31524
rect 26712 31210 26740 41262
rect 26896 41154 26924 41262
rect 27038 41200 27150 42000
rect 27682 41200 27794 42000
rect 28326 41200 28438 42000
rect 28970 41200 29082 42000
rect 30258 41200 30370 42000
rect 30902 41200 31014 42000
rect 31546 41200 31658 42000
rect 32190 41200 32302 42000
rect 32834 41200 32946 42000
rect 33478 41200 33590 42000
rect 34122 41200 34234 42000
rect 34766 41200 34878 42000
rect 35410 41200 35522 42000
rect 27080 41154 27108 41200
rect 26896 41126 27108 41154
rect 28264 38344 28316 38350
rect 28264 38286 28316 38292
rect 28276 37874 28304 38286
rect 28264 37868 28316 37874
rect 28264 37810 28316 37816
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 27816 35086 27844 36722
rect 27896 36168 27948 36174
rect 27896 36110 27948 36116
rect 27908 35698 27936 36110
rect 28368 35894 28396 41200
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 28460 37874 28488 38694
rect 28632 38208 28684 38214
rect 28632 38150 28684 38156
rect 28644 37942 28672 38150
rect 28632 37936 28684 37942
rect 28632 37878 28684 37884
rect 28448 37868 28500 37874
rect 28448 37810 28500 37816
rect 29012 37806 29040 41200
rect 31758 40896 31814 40905
rect 31758 40831 31814 40840
rect 31772 40118 31800 40831
rect 29736 40112 29788 40118
rect 29736 40054 29788 40060
rect 31760 40112 31812 40118
rect 31760 40054 31812 40060
rect 29000 37800 29052 37806
rect 29000 37742 29052 37748
rect 28368 35866 28488 35894
rect 27896 35692 27948 35698
rect 27896 35634 27948 35640
rect 28080 35624 28132 35630
rect 28080 35566 28132 35572
rect 28092 35290 28120 35566
rect 28080 35284 28132 35290
rect 28080 35226 28132 35232
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 27632 33522 27660 33934
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27816 33114 27844 33390
rect 27804 33108 27856 33114
rect 27804 33050 27856 33056
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26988 31346 27016 31758
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 26700 31204 26752 31210
rect 26700 31146 26752 31152
rect 26294 30492 26602 30501
rect 26294 30490 26300 30492
rect 26356 30490 26380 30492
rect 26436 30490 26460 30492
rect 26516 30490 26540 30492
rect 26596 30490 26602 30492
rect 26356 30438 26358 30490
rect 26538 30438 26540 30490
rect 26294 30436 26300 30438
rect 26356 30436 26380 30438
rect 26436 30436 26460 30438
rect 26516 30436 26540 30438
rect 26596 30436 26602 30438
rect 26294 30427 26602 30436
rect 27804 30388 27856 30394
rect 27804 30330 27856 30336
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 25412 29708 25464 29714
rect 25412 29650 25464 29656
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25240 29170 25268 29582
rect 25412 29572 25464 29578
rect 25412 29514 25464 29520
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25424 28762 25452 29514
rect 26294 29404 26602 29413
rect 26294 29402 26300 29404
rect 26356 29402 26380 29404
rect 26436 29402 26460 29404
rect 26516 29402 26540 29404
rect 26596 29402 26602 29404
rect 26356 29350 26358 29402
rect 26538 29350 26540 29402
rect 26294 29348 26300 29350
rect 26356 29348 26380 29350
rect 26436 29348 26460 29350
rect 26516 29348 26540 29350
rect 26596 29348 26602 29350
rect 26294 29339 26602 29348
rect 27080 29170 27108 29990
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27264 29238 27292 29446
rect 27252 29232 27304 29238
rect 27252 29174 27304 29180
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 25504 28960 25556 28966
rect 25504 28902 25556 28908
rect 25412 28756 25464 28762
rect 25412 28698 25464 28704
rect 25516 28626 25544 28902
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 27816 28558 27844 30330
rect 28460 29102 28488 35866
rect 29748 35766 29776 40054
rect 30518 39740 30826 39749
rect 30518 39738 30524 39740
rect 30580 39738 30604 39740
rect 30660 39738 30684 39740
rect 30740 39738 30764 39740
rect 30820 39738 30826 39740
rect 30580 39686 30582 39738
rect 30762 39686 30764 39738
rect 30518 39684 30524 39686
rect 30580 39684 30604 39686
rect 30660 39684 30684 39686
rect 30740 39684 30764 39686
rect 30820 39684 30826 39686
rect 30518 39675 30826 39684
rect 32876 39658 32904 41200
rect 31864 39630 32904 39658
rect 31758 38856 31814 38865
rect 31758 38791 31760 38800
rect 31812 38791 31814 38800
rect 31760 38762 31812 38768
rect 30518 38652 30826 38661
rect 30518 38650 30524 38652
rect 30580 38650 30604 38652
rect 30660 38650 30684 38652
rect 30740 38650 30764 38652
rect 30820 38650 30826 38652
rect 30580 38598 30582 38650
rect 30762 38598 30764 38650
rect 30518 38596 30524 38598
rect 30580 38596 30604 38598
rect 30660 38596 30684 38598
rect 30740 38596 30764 38598
rect 30820 38596 30826 38598
rect 30518 38587 30826 38596
rect 30288 38344 30340 38350
rect 30288 38286 30340 38292
rect 30300 37330 30328 38286
rect 30518 37564 30826 37573
rect 30518 37562 30524 37564
rect 30580 37562 30604 37564
rect 30660 37562 30684 37564
rect 30740 37562 30764 37564
rect 30820 37562 30826 37564
rect 30580 37510 30582 37562
rect 30762 37510 30764 37562
rect 30518 37508 30524 37510
rect 30580 37508 30604 37510
rect 30660 37508 30684 37510
rect 30740 37508 30764 37510
rect 30820 37508 30826 37510
rect 30518 37499 30826 37508
rect 30288 37324 30340 37330
rect 30288 37266 30340 37272
rect 29736 35760 29788 35766
rect 29736 35702 29788 35708
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 28448 29096 28500 29102
rect 28448 29038 28500 29044
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 27804 28552 27856 28558
rect 27804 28494 27856 28500
rect 25504 28484 25556 28490
rect 25504 28426 25556 28432
rect 25516 28218 25544 28426
rect 26294 28316 26602 28325
rect 26294 28314 26300 28316
rect 26356 28314 26380 28316
rect 26436 28314 26460 28316
rect 26516 28314 26540 28316
rect 26596 28314 26602 28316
rect 26356 28262 26358 28314
rect 26538 28262 26540 28314
rect 26294 28260 26300 28262
rect 26356 28260 26380 28262
rect 26436 28260 26460 28262
rect 26516 28260 26540 28262
rect 26596 28260 26602 28262
rect 26294 28251 26602 28260
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25412 28076 25464 28082
rect 25412 28018 25464 28024
rect 25424 24818 25452 28018
rect 26294 27228 26602 27237
rect 26294 27226 26300 27228
rect 26356 27226 26380 27228
rect 26436 27226 26460 27228
rect 26516 27226 26540 27228
rect 26596 27226 26602 27228
rect 26356 27174 26358 27226
rect 26538 27174 26540 27226
rect 26294 27172 26300 27174
rect 26356 27172 26380 27174
rect 26436 27172 26460 27174
rect 26516 27172 26540 27174
rect 26596 27172 26602 27174
rect 26294 27163 26602 27172
rect 26294 26140 26602 26149
rect 26294 26138 26300 26140
rect 26356 26138 26380 26140
rect 26436 26138 26460 26140
rect 26516 26138 26540 26140
rect 26596 26138 26602 26140
rect 26356 26086 26358 26138
rect 26538 26086 26540 26138
rect 26294 26084 26300 26086
rect 26356 26084 26380 26086
rect 26436 26084 26460 26086
rect 26516 26084 26540 26086
rect 26596 26084 26602 26086
rect 26294 26075 26602 26084
rect 26294 25052 26602 25061
rect 26294 25050 26300 25052
rect 26356 25050 26380 25052
rect 26436 25050 26460 25052
rect 26516 25050 26540 25052
rect 26596 25050 26602 25052
rect 26356 24998 26358 25050
rect 26538 24998 26540 25050
rect 26294 24996 26300 24998
rect 26356 24996 26380 24998
rect 26436 24996 26460 24998
rect 26516 24996 26540 24998
rect 26596 24996 26602 24998
rect 26294 24987 26602 24996
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 26294 23964 26602 23973
rect 26294 23962 26300 23964
rect 26356 23962 26380 23964
rect 26436 23962 26460 23964
rect 26516 23962 26540 23964
rect 26596 23962 26602 23964
rect 26356 23910 26358 23962
rect 26538 23910 26540 23962
rect 26294 23908 26300 23910
rect 26356 23908 26380 23910
rect 26436 23908 26460 23910
rect 26516 23908 26540 23910
rect 26596 23908 26602 23910
rect 26294 23899 26602 23908
rect 26294 22876 26602 22885
rect 26294 22874 26300 22876
rect 26356 22874 26380 22876
rect 26436 22874 26460 22876
rect 26516 22874 26540 22876
rect 26596 22874 26602 22876
rect 26356 22822 26358 22874
rect 26538 22822 26540 22874
rect 26294 22820 26300 22822
rect 26356 22820 26380 22822
rect 26436 22820 26460 22822
rect 26516 22820 26540 22822
rect 26596 22820 26602 22822
rect 26294 22811 26602 22820
rect 26294 21788 26602 21797
rect 26294 21786 26300 21788
rect 26356 21786 26380 21788
rect 26436 21786 26460 21788
rect 26516 21786 26540 21788
rect 26596 21786 26602 21788
rect 26356 21734 26358 21786
rect 26538 21734 26540 21786
rect 26294 21732 26300 21734
rect 26356 21732 26380 21734
rect 26436 21732 26460 21734
rect 26516 21732 26540 21734
rect 26596 21732 26602 21734
rect 26294 21723 26602 21732
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 22070 21244 22378 21253
rect 22070 21242 22076 21244
rect 22132 21242 22156 21244
rect 22212 21242 22236 21244
rect 22292 21242 22316 21244
rect 22372 21242 22378 21244
rect 22132 21190 22134 21242
rect 22314 21190 22316 21242
rect 22070 21188 22076 21190
rect 22132 21188 22156 21190
rect 22212 21188 22236 21190
rect 22292 21188 22316 21190
rect 22372 21188 22378 21190
rect 22070 21179 22378 21188
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20732 12458 20760 20402
rect 22070 20156 22378 20165
rect 22070 20154 22076 20156
rect 22132 20154 22156 20156
rect 22212 20154 22236 20156
rect 22292 20154 22316 20156
rect 22372 20154 22378 20156
rect 22132 20102 22134 20154
rect 22314 20102 22316 20154
rect 22070 20100 22076 20102
rect 22132 20100 22156 20102
rect 22212 20100 22236 20102
rect 22292 20100 22316 20102
rect 22372 20100 22378 20102
rect 22070 20091 22378 20100
rect 23492 19378 23520 21422
rect 26294 20700 26602 20709
rect 26294 20698 26300 20700
rect 26356 20698 26380 20700
rect 26436 20698 26460 20700
rect 26516 20698 26540 20700
rect 26596 20698 26602 20700
rect 26356 20646 26358 20698
rect 26538 20646 26540 20698
rect 26294 20644 26300 20646
rect 26356 20644 26380 20646
rect 26436 20644 26460 20646
rect 26516 20644 26540 20646
rect 26596 20644 26602 20646
rect 26294 20635 26602 20644
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24596 19922 24624 20198
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 24320 19514 24348 19722
rect 26294 19612 26602 19621
rect 26294 19610 26300 19612
rect 26356 19610 26380 19612
rect 26436 19610 26460 19612
rect 26516 19610 26540 19612
rect 26596 19610 26602 19612
rect 26356 19558 26358 19610
rect 26538 19558 26540 19610
rect 26294 19556 26300 19558
rect 26356 19556 26380 19558
rect 26436 19556 26460 19558
rect 26516 19556 26540 19558
rect 26596 19556 26602 19558
rect 26294 19547 26602 19556
rect 24308 19508 24360 19514
rect 24308 19450 24360 19456
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 22070 19068 22378 19077
rect 22070 19066 22076 19068
rect 22132 19066 22156 19068
rect 22212 19066 22236 19068
rect 22292 19066 22316 19068
rect 22372 19066 22378 19068
rect 22132 19014 22134 19066
rect 22314 19014 22316 19066
rect 22070 19012 22076 19014
rect 22132 19012 22156 19014
rect 22212 19012 22236 19014
rect 22292 19012 22316 19014
rect 22372 19012 22378 19014
rect 22070 19003 22378 19012
rect 26294 18524 26602 18533
rect 26294 18522 26300 18524
rect 26356 18522 26380 18524
rect 26436 18522 26460 18524
rect 26516 18522 26540 18524
rect 26596 18522 26602 18524
rect 26356 18470 26358 18522
rect 26538 18470 26540 18522
rect 26294 18468 26300 18470
rect 26356 18468 26380 18470
rect 26436 18468 26460 18470
rect 26516 18468 26540 18470
rect 26596 18468 26602 18470
rect 26294 18459 26602 18468
rect 22070 17980 22378 17989
rect 22070 17978 22076 17980
rect 22132 17978 22156 17980
rect 22212 17978 22236 17980
rect 22292 17978 22316 17980
rect 22372 17978 22378 17980
rect 22132 17926 22134 17978
rect 22314 17926 22316 17978
rect 22070 17924 22076 17926
rect 22132 17924 22156 17926
rect 22212 17924 22236 17926
rect 22292 17924 22316 17926
rect 22372 17924 22378 17926
rect 22070 17915 22378 17924
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 22070 16892 22378 16901
rect 22070 16890 22076 16892
rect 22132 16890 22156 16892
rect 22212 16890 22236 16892
rect 22292 16890 22316 16892
rect 22372 16890 22378 16892
rect 22132 16838 22134 16890
rect 22314 16838 22316 16890
rect 22070 16836 22076 16838
rect 22132 16836 22156 16838
rect 22212 16836 22236 16838
rect 22292 16836 22316 16838
rect 22372 16836 22378 16838
rect 22070 16827 22378 16836
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20824 15706 20852 15914
rect 22070 15804 22378 15813
rect 22070 15802 22076 15804
rect 22132 15802 22156 15804
rect 22212 15802 22236 15804
rect 22292 15802 22316 15804
rect 22372 15802 22378 15804
rect 22132 15750 22134 15802
rect 22314 15750 22316 15802
rect 22070 15748 22076 15750
rect 22132 15748 22156 15750
rect 22212 15748 22236 15750
rect 22292 15748 22316 15750
rect 22372 15748 22378 15750
rect 22070 15739 22378 15748
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20732 12430 20852 12458
rect 20824 11762 20852 12430
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10674 20760 11086
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17144 5234 17172 6326
rect 19720 5710 19748 6734
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 17846 5468 18154 5477
rect 17846 5466 17852 5468
rect 17908 5466 17932 5468
rect 17988 5466 18012 5468
rect 18068 5466 18092 5468
rect 18148 5466 18154 5468
rect 17908 5414 17910 5466
rect 18090 5414 18092 5466
rect 17846 5412 17852 5414
rect 17908 5412 17932 5414
rect 17988 5412 18012 5414
rect 18068 5412 18092 5414
rect 18148 5412 18154 5414
rect 17846 5403 18154 5412
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17846 4380 18154 4389
rect 17846 4378 17852 4380
rect 17908 4378 17932 4380
rect 17988 4378 18012 4380
rect 18068 4378 18092 4380
rect 18148 4378 18154 4380
rect 17908 4326 17910 4378
rect 18090 4326 18092 4378
rect 17846 4324 17852 4326
rect 17908 4324 17932 4326
rect 17988 4324 18012 4326
rect 18068 4324 18092 4326
rect 18148 4324 18154 4326
rect 17846 4315 18154 4324
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17604 3058 17632 3470
rect 17846 3292 18154 3301
rect 17846 3290 17852 3292
rect 17908 3290 17932 3292
rect 17988 3290 18012 3292
rect 18068 3290 18092 3292
rect 18148 3290 18154 3292
rect 17908 3238 17910 3290
rect 18090 3238 18092 3290
rect 17846 3236 17852 3238
rect 17908 3236 17932 3238
rect 17988 3236 18012 3238
rect 18068 3236 18092 3238
rect 18148 3236 18154 3238
rect 17846 3227 18154 3236
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 16960 2446 16988 2994
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16868 2230 17448 2258
rect 17420 800 17448 2230
rect 17846 2204 18154 2213
rect 17846 2202 17852 2204
rect 17908 2202 17932 2204
rect 17988 2202 18012 2204
rect 18068 2202 18092 2204
rect 18148 2202 18154 2204
rect 17908 2150 17910 2202
rect 18090 2150 18092 2202
rect 17846 2148 17852 2150
rect 17908 2148 17932 2150
rect 17988 2148 18012 2150
rect 18068 2148 18092 2150
rect 18148 2148 18154 2150
rect 17846 2139 18154 2148
rect 19996 800 20024 9454
rect 20824 9042 20852 11698
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11218 20944 11494
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 21008 7410 21036 15438
rect 22070 14716 22378 14725
rect 22070 14714 22076 14716
rect 22132 14714 22156 14716
rect 22212 14714 22236 14716
rect 22292 14714 22316 14716
rect 22372 14714 22378 14716
rect 22132 14662 22134 14714
rect 22314 14662 22316 14714
rect 22070 14660 22076 14662
rect 22132 14660 22156 14662
rect 22212 14660 22236 14662
rect 22292 14660 22316 14662
rect 22372 14660 22378 14662
rect 22070 14651 22378 14660
rect 22070 13628 22378 13637
rect 22070 13626 22076 13628
rect 22132 13626 22156 13628
rect 22212 13626 22236 13628
rect 22292 13626 22316 13628
rect 22372 13626 22378 13628
rect 22132 13574 22134 13626
rect 22314 13574 22316 13626
rect 22070 13572 22076 13574
rect 22132 13572 22156 13574
rect 22212 13572 22236 13574
rect 22292 13572 22316 13574
rect 22372 13572 22378 13574
rect 22070 13563 22378 13572
rect 25240 12866 25268 17478
rect 26294 17436 26602 17445
rect 26294 17434 26300 17436
rect 26356 17434 26380 17436
rect 26436 17434 26460 17436
rect 26516 17434 26540 17436
rect 26596 17434 26602 17436
rect 26356 17382 26358 17434
rect 26538 17382 26540 17434
rect 26294 17380 26300 17382
rect 26356 17380 26380 17382
rect 26436 17380 26460 17382
rect 26516 17380 26540 17382
rect 26596 17380 26602 17382
rect 26294 17371 26602 17380
rect 26294 16348 26602 16357
rect 26294 16346 26300 16348
rect 26356 16346 26380 16348
rect 26436 16346 26460 16348
rect 26516 16346 26540 16348
rect 26596 16346 26602 16348
rect 26356 16294 26358 16346
rect 26538 16294 26540 16346
rect 26294 16292 26300 16294
rect 26356 16292 26380 16294
rect 26436 16292 26460 16294
rect 26516 16292 26540 16294
rect 26596 16292 26602 16294
rect 26294 16283 26602 16292
rect 26294 15260 26602 15269
rect 26294 15258 26300 15260
rect 26356 15258 26380 15260
rect 26436 15258 26460 15260
rect 26516 15258 26540 15260
rect 26596 15258 26602 15260
rect 26356 15206 26358 15258
rect 26538 15206 26540 15258
rect 26294 15204 26300 15206
rect 26356 15204 26380 15206
rect 26436 15204 26460 15206
rect 26516 15204 26540 15206
rect 26596 15204 26602 15206
rect 26294 15195 26602 15204
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25516 14482 25544 14758
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25332 13938 25360 14350
rect 26294 14172 26602 14181
rect 26294 14170 26300 14172
rect 26356 14170 26380 14172
rect 26436 14170 26460 14172
rect 26516 14170 26540 14172
rect 26596 14170 26602 14172
rect 26356 14118 26358 14170
rect 26538 14118 26540 14170
rect 26294 14116 26300 14118
rect 26356 14116 26380 14118
rect 26436 14116 26460 14118
rect 26516 14116 26540 14118
rect 26596 14116 26602 14118
rect 26294 14107 26602 14116
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25976 13394 26004 13670
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 12986 25636 13194
rect 26294 13084 26602 13093
rect 26294 13082 26300 13084
rect 26356 13082 26380 13084
rect 26436 13082 26460 13084
rect 26516 13082 26540 13084
rect 26596 13082 26602 13084
rect 26356 13030 26358 13082
rect 26538 13030 26540 13082
rect 26294 13028 26300 13030
rect 26356 13028 26380 13030
rect 26436 13028 26460 13030
rect 26516 13028 26540 13030
rect 26596 13028 26602 13030
rect 26294 13019 26602 13028
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25240 12850 25360 12866
rect 25240 12844 25372 12850
rect 25240 12838 25320 12844
rect 25320 12786 25372 12792
rect 22070 12540 22378 12549
rect 22070 12538 22076 12540
rect 22132 12538 22156 12540
rect 22212 12538 22236 12540
rect 22292 12538 22316 12540
rect 22372 12538 22378 12540
rect 22132 12486 22134 12538
rect 22314 12486 22316 12538
rect 22070 12484 22076 12486
rect 22132 12484 22156 12486
rect 22212 12484 22236 12486
rect 22292 12484 22316 12486
rect 22372 12484 22378 12486
rect 22070 12475 22378 12484
rect 22070 11452 22378 11461
rect 22070 11450 22076 11452
rect 22132 11450 22156 11452
rect 22212 11450 22236 11452
rect 22292 11450 22316 11452
rect 22372 11450 22378 11452
rect 22132 11398 22134 11450
rect 22314 11398 22316 11450
rect 22070 11396 22076 11398
rect 22132 11396 22156 11398
rect 22212 11396 22236 11398
rect 22292 11396 22316 11398
rect 22372 11396 22378 11398
rect 22070 11387 22378 11396
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20088 6866 20116 7142
rect 20824 6866 20852 7142
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20640 800 20668 6666
rect 21284 870 21496 898
rect 21284 800 21312 870
rect 9876 734 10088 762
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21468 762 21496 870
rect 21744 762 21772 11154
rect 22070 10364 22378 10373
rect 22070 10362 22076 10364
rect 22132 10362 22156 10364
rect 22212 10362 22236 10364
rect 22292 10362 22316 10364
rect 22372 10362 22378 10364
rect 22132 10310 22134 10362
rect 22314 10310 22316 10362
rect 22070 10308 22076 10310
rect 22132 10308 22156 10310
rect 22212 10308 22236 10310
rect 22292 10308 22316 10310
rect 22372 10308 22378 10310
rect 22070 10299 22378 10308
rect 22070 9276 22378 9285
rect 22070 9274 22076 9276
rect 22132 9274 22156 9276
rect 22212 9274 22236 9276
rect 22292 9274 22316 9276
rect 22372 9274 22378 9276
rect 22132 9222 22134 9274
rect 22314 9222 22316 9274
rect 22070 9220 22076 9222
rect 22132 9220 22156 9222
rect 22212 9220 22236 9222
rect 22292 9220 22316 9222
rect 22372 9220 22378 9222
rect 22070 9211 22378 9220
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23952 8498 23980 8910
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24136 8566 24164 8774
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 22070 8188 22378 8197
rect 22070 8186 22076 8188
rect 22132 8186 22156 8188
rect 22212 8186 22236 8188
rect 22292 8186 22316 8188
rect 22372 8186 22378 8188
rect 22132 8134 22134 8186
rect 22314 8134 22316 8186
rect 22070 8132 22076 8134
rect 22132 8132 22156 8134
rect 22212 8132 22236 8134
rect 22292 8132 22316 8134
rect 22372 8132 22378 8134
rect 22070 8123 22378 8132
rect 22070 7100 22378 7109
rect 22070 7098 22076 7100
rect 22132 7098 22156 7100
rect 22212 7098 22236 7100
rect 22292 7098 22316 7100
rect 22372 7098 22378 7100
rect 22132 7046 22134 7098
rect 22314 7046 22316 7098
rect 22070 7044 22076 7046
rect 22132 7044 22156 7046
rect 22212 7044 22236 7046
rect 22292 7044 22316 7046
rect 22372 7044 22378 7046
rect 22070 7035 22378 7044
rect 22070 6012 22378 6021
rect 22070 6010 22076 6012
rect 22132 6010 22156 6012
rect 22212 6010 22236 6012
rect 22292 6010 22316 6012
rect 22372 6010 22378 6012
rect 22132 5958 22134 6010
rect 22314 5958 22316 6010
rect 22070 5956 22076 5958
rect 22132 5956 22156 5958
rect 22212 5956 22236 5958
rect 22292 5956 22316 5958
rect 22372 5956 22378 5958
rect 22070 5947 22378 5956
rect 22070 4924 22378 4933
rect 22070 4922 22076 4924
rect 22132 4922 22156 4924
rect 22212 4922 22236 4924
rect 22292 4922 22316 4924
rect 22372 4922 22378 4924
rect 22132 4870 22134 4922
rect 22314 4870 22316 4922
rect 22070 4868 22076 4870
rect 22132 4868 22156 4870
rect 22212 4868 22236 4870
rect 22292 4868 22316 4870
rect 22372 4868 22378 4870
rect 22070 4859 22378 4868
rect 22070 3836 22378 3845
rect 22070 3834 22076 3836
rect 22132 3834 22156 3836
rect 22212 3834 22236 3836
rect 22292 3834 22316 3836
rect 22372 3834 22378 3836
rect 22132 3782 22134 3834
rect 22314 3782 22316 3834
rect 22070 3780 22076 3782
rect 22132 3780 22156 3782
rect 22212 3780 22236 3782
rect 22292 3780 22316 3782
rect 22372 3780 22378 3782
rect 22070 3771 22378 3780
rect 22070 2748 22378 2757
rect 22070 2746 22076 2748
rect 22132 2746 22156 2748
rect 22212 2746 22236 2748
rect 22292 2746 22316 2748
rect 22372 2746 22378 2748
rect 22132 2694 22134 2746
rect 22314 2694 22316 2746
rect 22070 2692 22076 2694
rect 22132 2692 22156 2694
rect 22212 2692 22236 2694
rect 22292 2692 22316 2694
rect 22372 2692 22378 2694
rect 22070 2683 22378 2692
rect 24504 800 24532 8366
rect 25332 4622 25360 12786
rect 26294 11996 26602 12005
rect 26294 11994 26300 11996
rect 26356 11994 26380 11996
rect 26436 11994 26460 11996
rect 26516 11994 26540 11996
rect 26596 11994 26602 11996
rect 26356 11942 26358 11994
rect 26538 11942 26540 11994
rect 26294 11940 26300 11942
rect 26356 11940 26380 11942
rect 26436 11940 26460 11942
rect 26516 11940 26540 11942
rect 26596 11940 26602 11942
rect 26294 11931 26602 11940
rect 26294 10908 26602 10917
rect 26294 10906 26300 10908
rect 26356 10906 26380 10908
rect 26436 10906 26460 10908
rect 26516 10906 26540 10908
rect 26596 10906 26602 10908
rect 26356 10854 26358 10906
rect 26538 10854 26540 10906
rect 26294 10852 26300 10854
rect 26356 10852 26380 10854
rect 26436 10852 26460 10854
rect 26516 10852 26540 10854
rect 26596 10852 26602 10854
rect 26294 10843 26602 10852
rect 27080 10674 27108 24754
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27172 18290 27200 18702
rect 27344 18692 27396 18698
rect 27344 18634 27396 18640
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27172 17678 27200 18022
rect 27356 17882 27384 18634
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27816 17746 27844 28494
rect 29104 25906 29132 35022
rect 30300 32910 30328 37266
rect 31666 36816 31722 36825
rect 31666 36751 31722 36760
rect 30518 36476 30826 36485
rect 30518 36474 30524 36476
rect 30580 36474 30604 36476
rect 30660 36474 30684 36476
rect 30740 36474 30764 36476
rect 30820 36474 30826 36476
rect 30580 36422 30582 36474
rect 30762 36422 30764 36474
rect 30518 36420 30524 36422
rect 30580 36420 30604 36422
rect 30660 36420 30684 36422
rect 30740 36420 30764 36422
rect 30820 36420 30826 36422
rect 30518 36411 30826 36420
rect 30518 35388 30826 35397
rect 30518 35386 30524 35388
rect 30580 35386 30604 35388
rect 30660 35386 30684 35388
rect 30740 35386 30764 35388
rect 30820 35386 30826 35388
rect 30580 35334 30582 35386
rect 30762 35334 30764 35386
rect 30518 35332 30524 35334
rect 30580 35332 30604 35334
rect 30660 35332 30684 35334
rect 30740 35332 30764 35334
rect 30820 35332 30826 35334
rect 30518 35323 30826 35332
rect 31574 34776 31630 34785
rect 31574 34711 31630 34720
rect 30518 34300 30826 34309
rect 30518 34298 30524 34300
rect 30580 34298 30604 34300
rect 30660 34298 30684 34300
rect 30740 34298 30764 34300
rect 30820 34298 30826 34300
rect 30580 34246 30582 34298
rect 30762 34246 30764 34298
rect 30518 34244 30524 34246
rect 30580 34244 30604 34246
rect 30660 34244 30684 34246
rect 30740 34244 30764 34246
rect 30820 34244 30826 34246
rect 30518 34235 30826 34244
rect 30518 33212 30826 33221
rect 30518 33210 30524 33212
rect 30580 33210 30604 33212
rect 30660 33210 30684 33212
rect 30740 33210 30764 33212
rect 30820 33210 30826 33212
rect 30580 33158 30582 33210
rect 30762 33158 30764 33210
rect 30518 33156 30524 33158
rect 30580 33156 30604 33158
rect 30660 33156 30684 33158
rect 30740 33156 30764 33158
rect 30820 33156 30826 33158
rect 30518 33147 30826 33156
rect 29828 32904 29880 32910
rect 29828 32846 29880 32852
rect 30288 32904 30340 32910
rect 30288 32846 30340 32852
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29380 29170 29408 29582
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29552 29096 29604 29102
rect 29552 29038 29604 29044
rect 29564 28762 29592 29038
rect 29552 28756 29604 28762
rect 29552 28698 29604 28704
rect 29736 26376 29788 26382
rect 29736 26318 29788 26324
rect 29748 25906 29776 26318
rect 29092 25900 29144 25906
rect 29092 25842 29144 25848
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28368 20466 28396 20878
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 29104 20330 29132 25842
rect 29840 24206 29868 32846
rect 30518 32124 30826 32133
rect 30518 32122 30524 32124
rect 30580 32122 30604 32124
rect 30660 32122 30684 32124
rect 30740 32122 30764 32124
rect 30820 32122 30826 32124
rect 30580 32070 30582 32122
rect 30762 32070 30764 32122
rect 30518 32068 30524 32070
rect 30580 32068 30604 32070
rect 30660 32068 30684 32070
rect 30740 32068 30764 32070
rect 30820 32068 30826 32070
rect 30518 32059 30826 32068
rect 30518 31036 30826 31045
rect 30518 31034 30524 31036
rect 30580 31034 30604 31036
rect 30660 31034 30684 31036
rect 30740 31034 30764 31036
rect 30820 31034 30826 31036
rect 30580 30982 30582 31034
rect 30762 30982 30764 31034
rect 30518 30980 30524 30982
rect 30580 30980 30604 30982
rect 30660 30980 30684 30982
rect 30740 30980 30764 30982
rect 30820 30980 30826 30982
rect 30518 30971 30826 30980
rect 30518 29948 30826 29957
rect 30518 29946 30524 29948
rect 30580 29946 30604 29948
rect 30660 29946 30684 29948
rect 30740 29946 30764 29948
rect 30820 29946 30826 29948
rect 30580 29894 30582 29946
rect 30762 29894 30764 29946
rect 30518 29892 30524 29894
rect 30580 29892 30604 29894
rect 30660 29892 30684 29894
rect 30740 29892 30764 29894
rect 30820 29892 30826 29894
rect 30518 29883 30826 29892
rect 30518 28860 30826 28869
rect 30518 28858 30524 28860
rect 30580 28858 30604 28860
rect 30660 28858 30684 28860
rect 30740 28858 30764 28860
rect 30820 28858 30826 28860
rect 30580 28806 30582 28858
rect 30762 28806 30764 28858
rect 30518 28804 30524 28806
rect 30580 28804 30604 28806
rect 30660 28804 30684 28806
rect 30740 28804 30764 28806
rect 30820 28804 30826 28806
rect 30518 28795 30826 28804
rect 31588 28626 31616 34711
rect 31680 29238 31708 36751
rect 31864 32298 31892 39630
rect 32586 39536 32642 39545
rect 32586 39471 32642 39480
rect 32312 38344 32364 38350
rect 32312 38286 32364 38292
rect 32324 37874 32352 38286
rect 32312 37868 32364 37874
rect 32312 37810 32364 37816
rect 32496 37800 32548 37806
rect 32496 37742 32548 37748
rect 32508 37466 32536 37742
rect 32496 37460 32548 37466
rect 32496 37402 32548 37408
rect 32312 33448 32364 33454
rect 32310 33416 32312 33425
rect 32364 33416 32366 33425
rect 32310 33351 32366 33360
rect 32128 33312 32180 33318
rect 32128 33254 32180 33260
rect 32140 32978 32168 33254
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 31852 32292 31904 32298
rect 31852 32234 31904 32240
rect 32324 32026 32352 32302
rect 32312 32020 32364 32026
rect 32312 31962 32364 31968
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 31668 29232 31720 29238
rect 31668 29174 31720 29180
rect 31576 28620 31628 28626
rect 31576 28562 31628 28568
rect 30518 27772 30826 27781
rect 30518 27770 30524 27772
rect 30580 27770 30604 27772
rect 30660 27770 30684 27772
rect 30740 27770 30764 27772
rect 30820 27770 30826 27772
rect 30580 27718 30582 27770
rect 30762 27718 30764 27770
rect 30518 27716 30524 27718
rect 30580 27716 30604 27718
rect 30660 27716 30684 27718
rect 30740 27716 30764 27718
rect 30820 27716 30826 27718
rect 30518 27707 30826 27716
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 30518 26684 30826 26693
rect 30518 26682 30524 26684
rect 30580 26682 30604 26684
rect 30660 26682 30684 26684
rect 30740 26682 30764 26684
rect 30820 26682 30826 26684
rect 30580 26630 30582 26682
rect 30762 26630 30764 26682
rect 30518 26628 30524 26630
rect 30580 26628 30604 26630
rect 30660 26628 30684 26630
rect 30740 26628 30764 26630
rect 30820 26628 30826 26630
rect 30518 26619 30826 26628
rect 31312 26450 31340 26726
rect 31300 26444 31352 26450
rect 31300 26386 31352 26392
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 30518 25596 30826 25605
rect 30518 25594 30524 25596
rect 30580 25594 30604 25596
rect 30660 25594 30684 25596
rect 30740 25594 30764 25596
rect 30820 25594 30826 25596
rect 30580 25542 30582 25594
rect 30762 25542 30764 25594
rect 30518 25540 30524 25542
rect 30580 25540 30604 25542
rect 30660 25540 30684 25542
rect 30740 25540 30764 25542
rect 30820 25540 30826 25542
rect 30518 25531 30826 25540
rect 31758 25256 31814 25265
rect 31668 25220 31720 25226
rect 31758 25191 31814 25200
rect 31668 25162 31720 25168
rect 31680 24954 31708 25162
rect 31668 24948 31720 24954
rect 31668 24890 31720 24896
rect 31772 24834 31800 25191
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31680 24806 31800 24834
rect 30518 24508 30826 24517
rect 30518 24506 30524 24508
rect 30580 24506 30604 24508
rect 30660 24506 30684 24508
rect 30740 24506 30764 24508
rect 30820 24506 30826 24508
rect 30580 24454 30582 24506
rect 30762 24454 30764 24506
rect 30518 24452 30524 24454
rect 30580 24452 30604 24454
rect 30660 24452 30684 24454
rect 30740 24452 30764 24454
rect 30820 24452 30826 24454
rect 30518 24443 30826 24452
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29932 23798 29960 24006
rect 29920 23792 29972 23798
rect 29920 23734 29972 23740
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29184 23588 29236 23594
rect 29184 23530 29236 23536
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 27172 15026 27200 17614
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27724 17270 27752 17478
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27540 16794 27568 17070
rect 27528 16788 27580 16794
rect 27528 16730 27580 16736
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27816 10266 27844 10542
rect 27804 10260 27856 10266
rect 27804 10202 27856 10208
rect 28276 10062 28304 17614
rect 29196 16574 29224 23530
rect 29748 23322 29776 23598
rect 30518 23420 30826 23429
rect 30518 23418 30524 23420
rect 30580 23418 30604 23420
rect 30660 23418 30684 23420
rect 30740 23418 30764 23420
rect 30820 23418 30826 23420
rect 30580 23366 30582 23418
rect 30762 23366 30764 23418
rect 30518 23364 30524 23366
rect 30580 23364 30604 23366
rect 30660 23364 30684 23366
rect 30740 23364 30764 23366
rect 30820 23364 30826 23366
rect 30518 23355 30826 23364
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 30944 23254 30972 24142
rect 30932 23248 30984 23254
rect 30932 23190 30984 23196
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30852 22778 30880 22986
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 31128 22642 31156 24754
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 31116 22636 31168 22642
rect 31116 22578 31168 22584
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 19922 29592 20878
rect 29552 19916 29604 19922
rect 29552 19858 29604 19864
rect 30392 19446 30420 22578
rect 30518 22332 30826 22341
rect 30518 22330 30524 22332
rect 30580 22330 30604 22332
rect 30660 22330 30684 22332
rect 30740 22330 30764 22332
rect 30820 22330 30826 22332
rect 30580 22278 30582 22330
rect 30762 22278 30764 22330
rect 30518 22276 30524 22278
rect 30580 22276 30604 22278
rect 30660 22276 30684 22278
rect 30740 22276 30764 22278
rect 30820 22276 30826 22278
rect 30518 22267 30826 22276
rect 30518 21244 30826 21253
rect 30518 21242 30524 21244
rect 30580 21242 30604 21244
rect 30660 21242 30684 21244
rect 30740 21242 30764 21244
rect 30820 21242 30826 21244
rect 30580 21190 30582 21242
rect 30762 21190 30764 21242
rect 30518 21188 30524 21190
rect 30580 21188 30604 21190
rect 30660 21188 30684 21190
rect 30740 21188 30764 21190
rect 30820 21188 30826 21190
rect 30518 21179 30826 21188
rect 30518 20156 30826 20165
rect 30518 20154 30524 20156
rect 30580 20154 30604 20156
rect 30660 20154 30684 20156
rect 30740 20154 30764 20156
rect 30820 20154 30826 20156
rect 30580 20102 30582 20154
rect 30762 20102 30764 20154
rect 30518 20100 30524 20102
rect 30580 20100 30604 20102
rect 30660 20100 30684 20102
rect 30740 20100 30764 20102
rect 30820 20100 30826 20102
rect 30518 20091 30826 20100
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 30380 19440 30432 19446
rect 30380 19382 30432 19388
rect 29552 18080 29604 18086
rect 29552 18022 29604 18028
rect 29564 17746 29592 18022
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29196 16546 30236 16574
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 26294 9820 26602 9829
rect 26294 9818 26300 9820
rect 26356 9818 26380 9820
rect 26436 9818 26460 9820
rect 26516 9818 26540 9820
rect 26596 9818 26602 9820
rect 26356 9766 26358 9818
rect 26538 9766 26540 9818
rect 26294 9764 26300 9766
rect 26356 9764 26380 9766
rect 26436 9764 26460 9766
rect 26516 9764 26540 9766
rect 26596 9764 26602 9766
rect 26294 9755 26602 9764
rect 26294 8732 26602 8741
rect 26294 8730 26300 8732
rect 26356 8730 26380 8732
rect 26436 8730 26460 8732
rect 26516 8730 26540 8732
rect 26596 8730 26602 8732
rect 26356 8678 26358 8730
rect 26538 8678 26540 8730
rect 26294 8676 26300 8678
rect 26356 8676 26380 8678
rect 26436 8676 26460 8678
rect 26516 8676 26540 8678
rect 26596 8676 26602 8678
rect 26294 8667 26602 8676
rect 28276 8498 28304 9998
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29196 7818 29224 8230
rect 29748 7954 29776 8230
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 26294 7644 26602 7653
rect 26294 7642 26300 7644
rect 26356 7642 26380 7644
rect 26436 7642 26460 7644
rect 26516 7642 26540 7644
rect 26596 7642 26602 7644
rect 26356 7590 26358 7642
rect 26538 7590 26540 7642
rect 26294 7588 26300 7590
rect 26356 7588 26380 7590
rect 26436 7588 26460 7590
rect 26516 7588 26540 7590
rect 26596 7588 26602 7590
rect 26294 7579 26602 7588
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 26294 6556 26602 6565
rect 26294 6554 26300 6556
rect 26356 6554 26380 6556
rect 26436 6554 26460 6556
rect 26516 6554 26540 6556
rect 26596 6554 26602 6556
rect 26356 6502 26358 6554
rect 26538 6502 26540 6554
rect 26294 6500 26300 6502
rect 26356 6500 26380 6502
rect 26436 6500 26460 6502
rect 26516 6500 26540 6502
rect 26596 6500 26602 6502
rect 26294 6491 26602 6500
rect 27264 6322 27292 6734
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 29092 6248 29144 6254
rect 29092 6190 29144 6196
rect 26988 5914 27016 6190
rect 26976 5908 27028 5914
rect 26976 5850 27028 5856
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 26294 5468 26602 5477
rect 26294 5466 26300 5468
rect 26356 5466 26380 5468
rect 26436 5466 26460 5468
rect 26516 5466 26540 5468
rect 26596 5466 26602 5468
rect 26356 5414 26358 5466
rect 26538 5414 26540 5466
rect 26294 5412 26300 5414
rect 26356 5412 26380 5414
rect 26436 5412 26460 5414
rect 26516 5412 26540 5414
rect 26596 5412 26602 5414
rect 26294 5403 26602 5412
rect 27632 5370 27660 5646
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 27356 4826 27384 5102
rect 29104 5098 29132 6190
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 26294 4380 26602 4389
rect 26294 4378 26300 4380
rect 26356 4378 26380 4380
rect 26436 4378 26460 4380
rect 26516 4378 26540 4380
rect 26596 4378 26602 4380
rect 26356 4326 26358 4378
rect 26538 4326 26540 4378
rect 26294 4324 26300 4326
rect 26356 4324 26380 4326
rect 26436 4324 26460 4326
rect 26516 4324 26540 4326
rect 26596 4324 26602 4326
rect 26294 4315 26602 4324
rect 26294 3292 26602 3301
rect 26294 3290 26300 3292
rect 26356 3290 26380 3292
rect 26436 3290 26460 3292
rect 26516 3290 26540 3292
rect 26596 3290 26602 3292
rect 26356 3238 26358 3290
rect 26538 3238 26540 3290
rect 26294 3236 26300 3238
rect 26356 3236 26380 3238
rect 26436 3236 26460 3238
rect 26516 3236 26540 3238
rect 26596 3236 26602 3238
rect 26294 3227 26602 3236
rect 26294 2204 26602 2213
rect 26294 2202 26300 2204
rect 26356 2202 26380 2204
rect 26436 2202 26460 2204
rect 26516 2202 26540 2204
rect 26596 2202 26602 2204
rect 26356 2150 26358 2202
rect 26538 2150 26540 2202
rect 26294 2148 26300 2150
rect 26356 2148 26380 2150
rect 26436 2148 26460 2150
rect 26516 2148 26540 2150
rect 26596 2148 26602 2150
rect 26294 2139 26602 2148
rect 30208 2122 30236 16546
rect 30392 5234 30420 19382
rect 30518 19068 30826 19077
rect 30518 19066 30524 19068
rect 30580 19066 30604 19068
rect 30660 19066 30684 19068
rect 30740 19066 30764 19068
rect 30820 19066 30826 19068
rect 30580 19014 30582 19066
rect 30762 19014 30764 19066
rect 30518 19012 30524 19014
rect 30580 19012 30604 19014
rect 30660 19012 30684 19014
rect 30740 19012 30764 19014
rect 30820 19012 30826 19014
rect 30518 19003 30826 19012
rect 30518 17980 30826 17989
rect 30518 17978 30524 17980
rect 30580 17978 30604 17980
rect 30660 17978 30684 17980
rect 30740 17978 30764 17980
rect 30820 17978 30826 17980
rect 30580 17926 30582 17978
rect 30762 17926 30764 17978
rect 30518 17924 30524 17926
rect 30580 17924 30604 17926
rect 30660 17924 30684 17926
rect 30740 17924 30764 17926
rect 30820 17924 30826 17926
rect 30518 17915 30826 17924
rect 30518 16892 30826 16901
rect 30518 16890 30524 16892
rect 30580 16890 30604 16892
rect 30660 16890 30684 16892
rect 30740 16890 30764 16892
rect 30820 16890 30826 16892
rect 30580 16838 30582 16890
rect 30762 16838 30764 16890
rect 30518 16836 30524 16838
rect 30580 16836 30604 16838
rect 30660 16836 30684 16838
rect 30740 16836 30764 16838
rect 30820 16836 30826 16838
rect 30518 16827 30826 16836
rect 30518 15804 30826 15813
rect 30518 15802 30524 15804
rect 30580 15802 30604 15804
rect 30660 15802 30684 15804
rect 30740 15802 30764 15804
rect 30820 15802 30826 15804
rect 30580 15750 30582 15802
rect 30762 15750 30764 15802
rect 30518 15748 30524 15750
rect 30580 15748 30604 15750
rect 30660 15748 30684 15750
rect 30740 15748 30764 15750
rect 30820 15748 30826 15750
rect 30518 15739 30826 15748
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 30518 14716 30826 14725
rect 30518 14714 30524 14716
rect 30580 14714 30604 14716
rect 30660 14714 30684 14716
rect 30740 14714 30764 14716
rect 30820 14714 30826 14716
rect 30580 14662 30582 14714
rect 30762 14662 30764 14714
rect 30518 14660 30524 14662
rect 30580 14660 30604 14662
rect 30660 14660 30684 14662
rect 30740 14660 30764 14662
rect 30820 14660 30826 14662
rect 30518 14651 30826 14660
rect 30518 13628 30826 13637
rect 30518 13626 30524 13628
rect 30580 13626 30604 13628
rect 30660 13626 30684 13628
rect 30740 13626 30764 13628
rect 30820 13626 30826 13628
rect 30580 13574 30582 13626
rect 30762 13574 30764 13626
rect 30518 13572 30524 13574
rect 30580 13572 30604 13574
rect 30660 13572 30684 13574
rect 30740 13572 30764 13574
rect 30820 13572 30826 13574
rect 30518 13563 30826 13572
rect 30518 12540 30826 12549
rect 30518 12538 30524 12540
rect 30580 12538 30604 12540
rect 30660 12538 30684 12540
rect 30740 12538 30764 12540
rect 30820 12538 30826 12540
rect 30580 12486 30582 12538
rect 30762 12486 30764 12538
rect 30518 12484 30524 12486
rect 30580 12484 30604 12486
rect 30660 12484 30684 12486
rect 30740 12484 30764 12486
rect 30820 12484 30826 12486
rect 30518 12475 30826 12484
rect 30518 11452 30826 11461
rect 30518 11450 30524 11452
rect 30580 11450 30604 11452
rect 30660 11450 30684 11452
rect 30740 11450 30764 11452
rect 30820 11450 30826 11452
rect 30580 11398 30582 11450
rect 30762 11398 30764 11450
rect 30518 11396 30524 11398
rect 30580 11396 30604 11398
rect 30660 11396 30684 11398
rect 30740 11396 30764 11398
rect 30820 11396 30826 11398
rect 30518 11387 30826 11396
rect 30518 10364 30826 10373
rect 30518 10362 30524 10364
rect 30580 10362 30604 10364
rect 30660 10362 30684 10364
rect 30740 10362 30764 10364
rect 30820 10362 30826 10364
rect 30580 10310 30582 10362
rect 30762 10310 30764 10362
rect 30518 10308 30524 10310
rect 30580 10308 30604 10310
rect 30660 10308 30684 10310
rect 30740 10308 30764 10310
rect 30820 10308 30826 10310
rect 30518 10299 30826 10308
rect 30518 9276 30826 9285
rect 30518 9274 30524 9276
rect 30580 9274 30604 9276
rect 30660 9274 30684 9276
rect 30740 9274 30764 9276
rect 30820 9274 30826 9276
rect 30580 9222 30582 9274
rect 30762 9222 30764 9274
rect 30518 9220 30524 9222
rect 30580 9220 30604 9222
rect 30660 9220 30684 9222
rect 30740 9220 30764 9222
rect 30820 9220 30826 9222
rect 30518 9211 30826 9220
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30840 8900 30892 8906
rect 30840 8842 30892 8848
rect 30852 8634 30880 8842
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 30944 8498 30972 8910
rect 31036 8566 31064 14894
rect 31024 8560 31076 8566
rect 31024 8502 31076 8508
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30518 8188 30826 8197
rect 30518 8186 30524 8188
rect 30580 8186 30604 8188
rect 30660 8186 30684 8188
rect 30740 8186 30764 8188
rect 30820 8186 30826 8188
rect 30580 8134 30582 8186
rect 30762 8134 30764 8186
rect 30518 8132 30524 8134
rect 30580 8132 30604 8134
rect 30660 8132 30684 8134
rect 30740 8132 30764 8134
rect 30820 8132 30826 8134
rect 30518 8123 30826 8132
rect 30518 7100 30826 7109
rect 30518 7098 30524 7100
rect 30580 7098 30604 7100
rect 30660 7098 30684 7100
rect 30740 7098 30764 7100
rect 30820 7098 30826 7100
rect 30580 7046 30582 7098
rect 30762 7046 30764 7098
rect 30518 7044 30524 7046
rect 30580 7044 30604 7046
rect 30660 7044 30684 7046
rect 30740 7044 30764 7046
rect 30820 7044 30826 7046
rect 30518 7035 30826 7044
rect 31036 6914 31064 8502
rect 30944 6886 31064 6914
rect 30944 6798 30972 6886
rect 30932 6792 30984 6798
rect 30932 6734 30984 6740
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 30518 6012 30826 6021
rect 30518 6010 30524 6012
rect 30580 6010 30604 6012
rect 30660 6010 30684 6012
rect 30740 6010 30764 6012
rect 30820 6010 30826 6012
rect 30580 5958 30582 6010
rect 30762 5958 30764 6010
rect 30518 5956 30524 5958
rect 30580 5956 30604 5958
rect 30660 5956 30684 5958
rect 30740 5956 30764 5958
rect 30820 5956 30826 5958
rect 30518 5947 30826 5956
rect 30944 5778 30972 6598
rect 31220 5846 31248 6734
rect 31208 5840 31260 5846
rect 31208 5782 31260 5788
rect 30932 5772 30984 5778
rect 30932 5714 30984 5720
rect 30380 5228 30432 5234
rect 30380 5170 30432 5176
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30392 4758 30420 4966
rect 30518 4924 30826 4933
rect 30518 4922 30524 4924
rect 30580 4922 30604 4924
rect 30660 4922 30684 4924
rect 30740 4922 30764 4924
rect 30820 4922 30826 4924
rect 30580 4870 30582 4922
rect 30762 4870 30764 4922
rect 30518 4868 30524 4870
rect 30580 4868 30604 4870
rect 30660 4868 30684 4870
rect 30740 4868 30764 4870
rect 30820 4868 30826 4870
rect 30518 4859 30826 4868
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 30300 4146 30328 4558
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30518 3836 30826 3845
rect 30518 3834 30524 3836
rect 30580 3834 30604 3836
rect 30660 3834 30684 3836
rect 30740 3834 30764 3836
rect 30820 3834 30826 3836
rect 30580 3782 30582 3834
rect 30762 3782 30764 3834
rect 30518 3780 30524 3782
rect 30580 3780 30604 3782
rect 30660 3780 30684 3782
rect 30740 3780 30764 3782
rect 30820 3780 30826 3782
rect 30518 3771 30826 3780
rect 30518 2748 30826 2757
rect 30518 2746 30524 2748
rect 30580 2746 30604 2748
rect 30660 2746 30684 2748
rect 30740 2746 30764 2748
rect 30820 2746 30826 2748
rect 30580 2694 30582 2746
rect 30762 2694 30764 2746
rect 30518 2692 30524 2694
rect 30580 2692 30604 2694
rect 30660 2692 30684 2694
rect 30740 2692 30764 2694
rect 30820 2692 30826 2694
rect 30518 2683 30826 2692
rect 30208 2094 30328 2122
rect 30300 800 30328 2094
rect 30944 800 30972 4626
rect 21468 734 21772 762
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23174 0 23286 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 31404 785 31432 19722
rect 31680 18902 31708 24806
rect 31758 19816 31814 19825
rect 31758 19751 31814 19760
rect 31772 19718 31800 19751
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31668 18896 31720 18902
rect 31668 18838 31720 18844
rect 31956 14958 31984 25842
rect 32048 24206 32076 31758
rect 32312 30048 32364 30054
rect 32312 29990 32364 29996
rect 32324 29170 32352 29990
rect 32312 29164 32364 29170
rect 32312 29106 32364 29112
rect 32496 29096 32548 29102
rect 32496 29038 32548 29044
rect 32508 28218 32536 29038
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32220 26308 32272 26314
rect 32220 26250 32272 26256
rect 32232 26042 32260 26250
rect 32600 26234 32628 39471
rect 32954 34096 33010 34105
rect 32954 34031 33010 34040
rect 32416 26206 32628 26234
rect 32220 26036 32272 26042
rect 32220 25978 32272 25984
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 32048 23526 32076 24142
rect 32324 23730 32352 24550
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32036 23520 32088 23526
rect 32036 23462 32088 23468
rect 32048 18766 32076 23462
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32140 18290 32168 18702
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32324 18358 32352 18566
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 32312 17128 32364 17134
rect 32310 17096 32312 17105
rect 32364 17096 32366 17105
rect 32310 17031 32366 17040
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 16658 32352 16934
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32416 16046 32444 26206
rect 32968 25362 32996 34031
rect 33046 32056 33102 32065
rect 33046 31991 33102 32000
rect 33060 29714 33088 31991
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 33520 28626 33548 41200
rect 34164 38298 34192 41200
rect 34072 38270 34192 38298
rect 34072 38010 34100 38270
rect 34150 38176 34206 38185
rect 34150 38111 34206 38120
rect 34060 38004 34112 38010
rect 34060 37946 34112 37952
rect 34164 37942 34192 38111
rect 34152 37936 34204 37942
rect 34152 37878 34204 37884
rect 33692 32836 33744 32842
rect 33692 32778 33744 32784
rect 33704 32745 33732 32778
rect 33690 32736 33746 32745
rect 33690 32671 33746 32680
rect 34150 31376 34206 31385
rect 34150 31311 34206 31320
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 33784 30048 33836 30054
rect 33784 29990 33836 29996
rect 33796 28626 33824 29990
rect 33980 29714 34008 30670
rect 33968 29708 34020 29714
rect 33968 29650 34020 29656
rect 33968 29572 34020 29578
rect 33968 29514 34020 29520
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33784 28620 33836 28626
rect 33784 28562 33836 28568
rect 33416 28484 33468 28490
rect 33416 28426 33468 28432
rect 33428 28218 33456 28426
rect 33980 28218 34008 29514
rect 34164 29238 34192 31311
rect 34152 29232 34204 29238
rect 34152 29174 34204 29180
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 33140 28076 33192 28082
rect 33140 28018 33192 28024
rect 33324 28076 33376 28082
rect 33324 28018 33376 28024
rect 33046 27976 33102 27985
rect 33046 27911 33102 27920
rect 33060 26450 33088 27911
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33048 25968 33100 25974
rect 33046 25936 33048 25945
rect 33100 25936 33102 25945
rect 33046 25871 33102 25880
rect 32956 25356 33008 25362
rect 32956 25298 33008 25304
rect 32678 24576 32734 24585
rect 32678 24511 32734 24520
rect 32496 24064 32548 24070
rect 32496 24006 32548 24012
rect 32508 23798 32536 24006
rect 32496 23792 32548 23798
rect 32496 23734 32548 23740
rect 32692 23186 32720 24511
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32680 23180 32732 23186
rect 32680 23122 32732 23128
rect 32496 22976 32548 22982
rect 32496 22918 32548 22924
rect 32508 22710 32536 22918
rect 32496 22704 32548 22710
rect 32496 22646 32548 22652
rect 32784 22574 32812 24142
rect 33152 23118 33180 28018
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 32772 22568 32824 22574
rect 32772 22510 32824 22516
rect 32956 20528 33008 20534
rect 32954 20496 32956 20505
rect 33008 20496 33010 20505
rect 32954 20431 33010 20440
rect 33048 19304 33100 19310
rect 33048 19246 33100 19252
rect 33060 19145 33088 19246
rect 33046 19136 33102 19145
rect 33046 19071 33102 19080
rect 33046 17776 33102 17785
rect 33046 17711 33048 17720
rect 33100 17711 33102 17720
rect 33048 17682 33100 17688
rect 32772 16516 32824 16522
rect 32772 16458 32824 16464
rect 32784 16250 32812 16458
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 33152 16182 33180 23054
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33244 18970 33272 19246
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 33336 18766 33364 28018
rect 34150 23896 34206 23905
rect 34150 23831 34206 23840
rect 34164 23798 34192 23831
rect 34152 23792 34204 23798
rect 34152 23734 34204 23740
rect 34150 23216 34206 23225
rect 34150 23151 34206 23160
rect 34164 22710 34192 23151
rect 34152 22704 34204 22710
rect 34152 22646 34204 22652
rect 34152 19304 34204 19310
rect 34152 19246 34204 19252
rect 34164 18970 34192 19246
rect 34152 18964 34204 18970
rect 34152 18906 34204 18912
rect 33324 18760 33376 18766
rect 33324 18702 33376 18708
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 33140 16176 33192 16182
rect 33140 16118 33192 16124
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 31944 14952 31996 14958
rect 31944 14894 31996 14900
rect 31758 14376 31814 14385
rect 31758 14311 31760 14320
rect 31812 14311 31814 14320
rect 31760 14282 31812 14288
rect 32312 13728 32364 13734
rect 32312 13670 32364 13676
rect 32770 13696 32826 13705
rect 32324 12850 32352 13670
rect 32770 13631 32826 13640
rect 32784 13394 32812 13631
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 33048 13388 33100 13394
rect 33048 13330 33100 13336
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32508 12442 32536 12718
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 33060 12345 33088 13330
rect 33046 12336 33102 12345
rect 33046 12271 33102 12280
rect 33796 12238 33824 18702
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 31668 10600 31720 10606
rect 31668 10542 31720 10548
rect 31680 8922 31708 10542
rect 31758 8936 31814 8945
rect 31680 8894 31758 8922
rect 31758 8871 31814 8880
rect 32508 6746 32536 12174
rect 32772 8900 32824 8906
rect 32772 8842 32824 8848
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32692 6866 32720 7142
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 32416 6718 32536 6746
rect 32588 6724 32640 6730
rect 32416 6390 32444 6718
rect 32588 6666 32640 6672
rect 32600 6458 32628 6666
rect 32588 6452 32640 6458
rect 32588 6394 32640 6400
rect 32128 6384 32180 6390
rect 32128 6326 32180 6332
rect 32404 6384 32456 6390
rect 32404 6326 32456 6332
rect 32140 4146 32168 6326
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31772 2145 31800 2586
rect 31758 2136 31814 2145
rect 31758 2071 31814 2080
rect 32232 800 32260 5714
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32324 4865 32352 5102
rect 32404 5092 32456 5098
rect 32404 5034 32456 5040
rect 32310 4856 32366 4865
rect 32310 4791 32366 4800
rect 32416 4185 32444 5034
rect 32402 4176 32458 4185
rect 32402 4111 32458 4120
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32508 3602 32536 3878
rect 32496 3596 32548 3602
rect 32496 3538 32548 3544
rect 32784 3482 32812 8842
rect 33048 7812 33100 7818
rect 33048 7754 33100 7760
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 32876 3670 32904 3878
rect 32864 3664 32916 3670
rect 32864 3606 32916 3612
rect 33060 3505 33088 7754
rect 33888 6914 33916 18158
rect 34152 16516 34204 16522
rect 34152 16458 34204 16464
rect 34164 16425 34192 16458
rect 34150 16416 34206 16425
rect 34150 16351 34206 16360
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 33980 13394 34008 13670
rect 33968 13388 34020 13394
rect 33968 13330 34020 13336
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33980 12442 34008 13194
rect 34150 13016 34206 13025
rect 34150 12951 34206 12960
rect 34164 12918 34192 12951
rect 34152 12912 34204 12918
rect 34152 12854 34204 12860
rect 33968 12436 34020 12442
rect 33968 12378 34020 12384
rect 33888 6886 34008 6914
rect 33046 3496 33102 3505
rect 32784 3454 32904 3482
rect 32876 800 32904 3454
rect 33046 3431 33102 3440
rect 31390 776 31446 785
rect 31390 711 31446 720
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 33980 105 34008 6886
rect 34150 6896 34206 6905
rect 34150 6831 34152 6840
rect 34204 6831 34206 6840
rect 34152 6802 34204 6808
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 34808 800 34836 3402
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 35452 800 35480 2926
rect 33966 96 34022 105
rect 33966 31 34022 40
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
<< via2 >>
rect 3606 41520 3662 41576
rect 3330 37440 3386 37496
rect 1858 36100 1914 36136
rect 1858 36080 1860 36100
rect 1860 36080 1912 36100
rect 1912 36080 1914 36100
rect 3330 35400 3386 35456
rect 1858 14320 1914 14376
rect 2778 13640 2834 13696
rect 2778 10920 2834 10976
rect 1858 8880 1914 8936
rect 3422 34040 3478 34096
rect 3422 32000 3478 32056
rect 3422 31320 3478 31376
rect 3422 25200 3478 25256
rect 4066 40840 4122 40896
rect 5180 39738 5236 39740
rect 5260 39738 5316 39740
rect 5340 39738 5396 39740
rect 5420 39738 5476 39740
rect 5180 39686 5226 39738
rect 5226 39686 5236 39738
rect 5260 39686 5290 39738
rect 5290 39686 5302 39738
rect 5302 39686 5316 39738
rect 5340 39686 5354 39738
rect 5354 39686 5366 39738
rect 5366 39686 5396 39738
rect 5420 39686 5430 39738
rect 5430 39686 5476 39738
rect 5180 39684 5236 39686
rect 5260 39684 5316 39686
rect 5340 39684 5396 39686
rect 5420 39684 5476 39686
rect 5180 38650 5236 38652
rect 5260 38650 5316 38652
rect 5340 38650 5396 38652
rect 5420 38650 5476 38652
rect 5180 38598 5226 38650
rect 5226 38598 5236 38650
rect 5260 38598 5290 38650
rect 5290 38598 5302 38650
rect 5302 38598 5316 38650
rect 5340 38598 5354 38650
rect 5354 38598 5366 38650
rect 5366 38598 5396 38650
rect 5420 38598 5430 38650
rect 5430 38598 5476 38650
rect 5180 38596 5236 38598
rect 5260 38596 5316 38598
rect 5340 38596 5396 38598
rect 5420 38596 5476 38598
rect 5180 37562 5236 37564
rect 5260 37562 5316 37564
rect 5340 37562 5396 37564
rect 5420 37562 5476 37564
rect 5180 37510 5226 37562
rect 5226 37510 5236 37562
rect 5260 37510 5290 37562
rect 5290 37510 5302 37562
rect 5302 37510 5316 37562
rect 5340 37510 5354 37562
rect 5354 37510 5366 37562
rect 5366 37510 5396 37562
rect 5420 37510 5430 37562
rect 5430 37510 5476 37562
rect 5180 37508 5236 37510
rect 5260 37508 5316 37510
rect 5340 37508 5396 37510
rect 5420 37508 5476 37510
rect 4066 36760 4122 36816
rect 5180 36474 5236 36476
rect 5260 36474 5316 36476
rect 5340 36474 5396 36476
rect 5420 36474 5476 36476
rect 5180 36422 5226 36474
rect 5226 36422 5236 36474
rect 5260 36422 5290 36474
rect 5290 36422 5302 36474
rect 5302 36422 5316 36474
rect 5340 36422 5354 36474
rect 5354 36422 5366 36474
rect 5366 36422 5396 36474
rect 5420 36422 5430 36474
rect 5430 36422 5476 36474
rect 5180 36420 5236 36422
rect 5260 36420 5316 36422
rect 5340 36420 5396 36422
rect 5420 36420 5476 36422
rect 5180 35386 5236 35388
rect 5260 35386 5316 35388
rect 5340 35386 5396 35388
rect 5420 35386 5476 35388
rect 5180 35334 5226 35386
rect 5226 35334 5236 35386
rect 5260 35334 5290 35386
rect 5290 35334 5302 35386
rect 5302 35334 5316 35386
rect 5340 35334 5354 35386
rect 5354 35334 5366 35386
rect 5366 35334 5396 35386
rect 5420 35334 5430 35386
rect 5430 35334 5476 35386
rect 5180 35332 5236 35334
rect 5260 35332 5316 35334
rect 5340 35332 5396 35334
rect 5420 35332 5476 35334
rect 5180 34298 5236 34300
rect 5260 34298 5316 34300
rect 5340 34298 5396 34300
rect 5420 34298 5476 34300
rect 5180 34246 5226 34298
rect 5226 34246 5236 34298
rect 5260 34246 5290 34298
rect 5290 34246 5302 34298
rect 5302 34246 5316 34298
rect 5340 34246 5354 34298
rect 5354 34246 5366 34298
rect 5366 34246 5396 34298
rect 5420 34246 5430 34298
rect 5430 34246 5476 34298
rect 5180 34244 5236 34246
rect 5260 34244 5316 34246
rect 5340 34244 5396 34246
rect 5420 34244 5476 34246
rect 5180 33210 5236 33212
rect 5260 33210 5316 33212
rect 5340 33210 5396 33212
rect 5420 33210 5476 33212
rect 5180 33158 5226 33210
rect 5226 33158 5236 33210
rect 5260 33158 5290 33210
rect 5290 33158 5302 33210
rect 5302 33158 5316 33210
rect 5340 33158 5354 33210
rect 5354 33158 5366 33210
rect 5366 33158 5396 33210
rect 5420 33158 5430 33210
rect 5430 33158 5476 33210
rect 5180 33156 5236 33158
rect 5260 33156 5316 33158
rect 5340 33156 5396 33158
rect 5420 33156 5476 33158
rect 5180 32122 5236 32124
rect 5260 32122 5316 32124
rect 5340 32122 5396 32124
rect 5420 32122 5476 32124
rect 5180 32070 5226 32122
rect 5226 32070 5236 32122
rect 5260 32070 5290 32122
rect 5290 32070 5302 32122
rect 5302 32070 5316 32122
rect 5340 32070 5354 32122
rect 5354 32070 5366 32122
rect 5366 32070 5396 32122
rect 5420 32070 5430 32122
rect 5430 32070 5476 32122
rect 5180 32068 5236 32070
rect 5260 32068 5316 32070
rect 5340 32068 5396 32070
rect 5420 32068 5476 32070
rect 5180 31034 5236 31036
rect 5260 31034 5316 31036
rect 5340 31034 5396 31036
rect 5420 31034 5476 31036
rect 5180 30982 5226 31034
rect 5226 30982 5236 31034
rect 5260 30982 5290 31034
rect 5290 30982 5302 31034
rect 5302 30982 5316 31034
rect 5340 30982 5354 31034
rect 5354 30982 5366 31034
rect 5366 30982 5396 31034
rect 5420 30982 5430 31034
rect 5430 30982 5476 31034
rect 5180 30980 5236 30982
rect 5260 30980 5316 30982
rect 5340 30980 5396 30982
rect 5420 30980 5476 30982
rect 5180 29946 5236 29948
rect 5260 29946 5316 29948
rect 5340 29946 5396 29948
rect 5420 29946 5476 29948
rect 5180 29894 5226 29946
rect 5226 29894 5236 29946
rect 5260 29894 5290 29946
rect 5290 29894 5302 29946
rect 5302 29894 5316 29946
rect 5340 29894 5354 29946
rect 5354 29894 5366 29946
rect 5366 29894 5396 29946
rect 5420 29894 5430 29946
rect 5430 29894 5476 29946
rect 5180 29892 5236 29894
rect 5260 29892 5316 29894
rect 5340 29892 5396 29894
rect 5420 29892 5476 29894
rect 5180 28858 5236 28860
rect 5260 28858 5316 28860
rect 5340 28858 5396 28860
rect 5420 28858 5476 28860
rect 5180 28806 5226 28858
rect 5226 28806 5236 28858
rect 5260 28806 5290 28858
rect 5290 28806 5302 28858
rect 5302 28806 5316 28858
rect 5340 28806 5354 28858
rect 5354 28806 5366 28858
rect 5366 28806 5396 28858
rect 5420 28806 5430 28858
rect 5430 28806 5476 28858
rect 5180 28804 5236 28806
rect 5260 28804 5316 28806
rect 5340 28804 5396 28806
rect 5420 28804 5476 28806
rect 5180 27770 5236 27772
rect 5260 27770 5316 27772
rect 5340 27770 5396 27772
rect 5420 27770 5476 27772
rect 5180 27718 5226 27770
rect 5226 27718 5236 27770
rect 5260 27718 5290 27770
rect 5290 27718 5302 27770
rect 5302 27718 5316 27770
rect 5340 27718 5354 27770
rect 5354 27718 5366 27770
rect 5366 27718 5396 27770
rect 5420 27718 5430 27770
rect 5430 27718 5476 27770
rect 5180 27716 5236 27718
rect 5260 27716 5316 27718
rect 5340 27716 5396 27718
rect 5420 27716 5476 27718
rect 5180 26682 5236 26684
rect 5260 26682 5316 26684
rect 5340 26682 5396 26684
rect 5420 26682 5476 26684
rect 5180 26630 5226 26682
rect 5226 26630 5236 26682
rect 5260 26630 5290 26682
rect 5290 26630 5302 26682
rect 5302 26630 5316 26682
rect 5340 26630 5354 26682
rect 5354 26630 5366 26682
rect 5366 26630 5396 26682
rect 5420 26630 5430 26682
rect 5430 26630 5476 26682
rect 5180 26628 5236 26630
rect 5260 26628 5316 26630
rect 5340 26628 5396 26630
rect 5420 26628 5476 26630
rect 5180 25594 5236 25596
rect 5260 25594 5316 25596
rect 5340 25594 5396 25596
rect 5420 25594 5476 25596
rect 5180 25542 5226 25594
rect 5226 25542 5236 25594
rect 5260 25542 5290 25594
rect 5290 25542 5302 25594
rect 5302 25542 5316 25594
rect 5340 25542 5354 25594
rect 5354 25542 5366 25594
rect 5366 25542 5396 25594
rect 5420 25542 5430 25594
rect 5430 25542 5476 25594
rect 5180 25540 5236 25542
rect 5260 25540 5316 25542
rect 5340 25540 5396 25542
rect 5420 25540 5476 25542
rect 5180 24506 5236 24508
rect 5260 24506 5316 24508
rect 5340 24506 5396 24508
rect 5420 24506 5476 24508
rect 5180 24454 5226 24506
rect 5226 24454 5236 24506
rect 5260 24454 5290 24506
rect 5290 24454 5302 24506
rect 5302 24454 5316 24506
rect 5340 24454 5354 24506
rect 5354 24454 5366 24506
rect 5366 24454 5396 24506
rect 5420 24454 5430 24506
rect 5430 24454 5476 24506
rect 5180 24452 5236 24454
rect 5260 24452 5316 24454
rect 5340 24452 5396 24454
rect 5420 24452 5476 24454
rect 5180 23418 5236 23420
rect 5260 23418 5316 23420
rect 5340 23418 5396 23420
rect 5420 23418 5476 23420
rect 5180 23366 5226 23418
rect 5226 23366 5236 23418
rect 5260 23366 5290 23418
rect 5290 23366 5302 23418
rect 5302 23366 5316 23418
rect 5340 23366 5354 23418
rect 5354 23366 5366 23418
rect 5366 23366 5396 23418
rect 5420 23366 5430 23418
rect 5430 23366 5476 23418
rect 5180 23364 5236 23366
rect 5260 23364 5316 23366
rect 5340 23364 5396 23366
rect 5420 23364 5476 23366
rect 5180 22330 5236 22332
rect 5260 22330 5316 22332
rect 5340 22330 5396 22332
rect 5420 22330 5476 22332
rect 5180 22278 5226 22330
rect 5226 22278 5236 22330
rect 5260 22278 5290 22330
rect 5290 22278 5302 22330
rect 5302 22278 5316 22330
rect 5340 22278 5354 22330
rect 5354 22278 5366 22330
rect 5366 22278 5396 22330
rect 5420 22278 5430 22330
rect 5430 22278 5476 22330
rect 5180 22276 5236 22278
rect 5260 22276 5316 22278
rect 5340 22276 5396 22278
rect 5420 22276 5476 22278
rect 5180 21242 5236 21244
rect 5260 21242 5316 21244
rect 5340 21242 5396 21244
rect 5420 21242 5476 21244
rect 5180 21190 5226 21242
rect 5226 21190 5236 21242
rect 5260 21190 5290 21242
rect 5290 21190 5302 21242
rect 5302 21190 5316 21242
rect 5340 21190 5354 21242
rect 5354 21190 5366 21242
rect 5366 21190 5396 21242
rect 5420 21190 5430 21242
rect 5430 21190 5476 21242
rect 5180 21188 5236 21190
rect 5260 21188 5316 21190
rect 5340 21188 5396 21190
rect 5420 21188 5476 21190
rect 5180 20154 5236 20156
rect 5260 20154 5316 20156
rect 5340 20154 5396 20156
rect 5420 20154 5476 20156
rect 5180 20102 5226 20154
rect 5226 20102 5236 20154
rect 5260 20102 5290 20154
rect 5290 20102 5302 20154
rect 5302 20102 5316 20154
rect 5340 20102 5354 20154
rect 5354 20102 5366 20154
rect 5366 20102 5396 20154
rect 5420 20102 5430 20154
rect 5430 20102 5476 20154
rect 5180 20100 5236 20102
rect 5260 20100 5316 20102
rect 5340 20100 5396 20102
rect 5420 20100 5476 20102
rect 3422 19080 3478 19136
rect 5180 19066 5236 19068
rect 5260 19066 5316 19068
rect 5340 19066 5396 19068
rect 5420 19066 5476 19068
rect 5180 19014 5226 19066
rect 5226 19014 5236 19066
rect 5260 19014 5290 19066
rect 5290 19014 5302 19066
rect 5302 19014 5316 19066
rect 5340 19014 5354 19066
rect 5354 19014 5366 19066
rect 5366 19014 5396 19066
rect 5420 19014 5430 19066
rect 5430 19014 5476 19066
rect 5180 19012 5236 19014
rect 5260 19012 5316 19014
rect 5340 19012 5396 19014
rect 5420 19012 5476 19014
rect 3422 18400 3478 18456
rect 5180 17978 5236 17980
rect 5260 17978 5316 17980
rect 5340 17978 5396 17980
rect 5420 17978 5476 17980
rect 5180 17926 5226 17978
rect 5226 17926 5236 17978
rect 5260 17926 5290 17978
rect 5290 17926 5302 17978
rect 5302 17926 5316 17978
rect 5340 17926 5354 17978
rect 5354 17926 5366 17978
rect 5366 17926 5396 17978
rect 5420 17926 5430 17978
rect 5430 17926 5476 17978
rect 5180 17924 5236 17926
rect 5260 17924 5316 17926
rect 5340 17924 5396 17926
rect 5420 17924 5476 17926
rect 3238 17040 3294 17096
rect 5180 16890 5236 16892
rect 5260 16890 5316 16892
rect 5340 16890 5396 16892
rect 5420 16890 5476 16892
rect 5180 16838 5226 16890
rect 5226 16838 5236 16890
rect 5260 16838 5290 16890
rect 5290 16838 5302 16890
rect 5302 16838 5316 16890
rect 5340 16838 5354 16890
rect 5354 16838 5366 16890
rect 5366 16838 5396 16890
rect 5420 16838 5430 16890
rect 5430 16838 5476 16890
rect 5180 16836 5236 16838
rect 5260 16836 5316 16838
rect 5340 16836 5396 16838
rect 5420 16836 5476 16838
rect 4066 15680 4122 15736
rect 5180 15802 5236 15804
rect 5260 15802 5316 15804
rect 5340 15802 5396 15804
rect 5420 15802 5476 15804
rect 5180 15750 5226 15802
rect 5226 15750 5236 15802
rect 5260 15750 5290 15802
rect 5290 15750 5302 15802
rect 5302 15750 5316 15802
rect 5340 15750 5354 15802
rect 5354 15750 5366 15802
rect 5366 15750 5396 15802
rect 5420 15750 5430 15802
rect 5430 15750 5476 15802
rect 5180 15748 5236 15750
rect 5260 15748 5316 15750
rect 5340 15748 5396 15750
rect 5420 15748 5476 15750
rect 5180 14714 5236 14716
rect 5260 14714 5316 14716
rect 5340 14714 5396 14716
rect 5420 14714 5476 14716
rect 5180 14662 5226 14714
rect 5226 14662 5236 14714
rect 5260 14662 5290 14714
rect 5290 14662 5302 14714
rect 5302 14662 5316 14714
rect 5340 14662 5354 14714
rect 5354 14662 5366 14714
rect 5366 14662 5396 14714
rect 5420 14662 5430 14714
rect 5430 14662 5476 14714
rect 5180 14660 5236 14662
rect 5260 14660 5316 14662
rect 5340 14660 5396 14662
rect 5420 14660 5476 14662
rect 5180 13626 5236 13628
rect 5260 13626 5316 13628
rect 5340 13626 5396 13628
rect 5420 13626 5476 13628
rect 5180 13574 5226 13626
rect 5226 13574 5236 13626
rect 5260 13574 5290 13626
rect 5290 13574 5302 13626
rect 5302 13574 5316 13626
rect 5340 13574 5354 13626
rect 5354 13574 5366 13626
rect 5366 13574 5396 13626
rect 5420 13574 5430 13626
rect 5430 13574 5476 13626
rect 5180 13572 5236 13574
rect 5260 13572 5316 13574
rect 5340 13572 5396 13574
rect 5420 13572 5476 13574
rect 13628 39738 13684 39740
rect 13708 39738 13764 39740
rect 13788 39738 13844 39740
rect 13868 39738 13924 39740
rect 13628 39686 13674 39738
rect 13674 39686 13684 39738
rect 13708 39686 13738 39738
rect 13738 39686 13750 39738
rect 13750 39686 13764 39738
rect 13788 39686 13802 39738
rect 13802 39686 13814 39738
rect 13814 39686 13844 39738
rect 13868 39686 13878 39738
rect 13878 39686 13924 39738
rect 13628 39684 13684 39686
rect 13708 39684 13764 39686
rect 13788 39684 13844 39686
rect 13868 39684 13924 39686
rect 9404 39194 9460 39196
rect 9484 39194 9540 39196
rect 9564 39194 9620 39196
rect 9644 39194 9700 39196
rect 9404 39142 9450 39194
rect 9450 39142 9460 39194
rect 9484 39142 9514 39194
rect 9514 39142 9526 39194
rect 9526 39142 9540 39194
rect 9564 39142 9578 39194
rect 9578 39142 9590 39194
rect 9590 39142 9620 39194
rect 9644 39142 9654 39194
rect 9654 39142 9700 39194
rect 9404 39140 9460 39142
rect 9484 39140 9540 39142
rect 9564 39140 9620 39142
rect 9644 39140 9700 39142
rect 13628 38650 13684 38652
rect 13708 38650 13764 38652
rect 13788 38650 13844 38652
rect 13868 38650 13924 38652
rect 13628 38598 13674 38650
rect 13674 38598 13684 38650
rect 13708 38598 13738 38650
rect 13738 38598 13750 38650
rect 13750 38598 13764 38650
rect 13788 38598 13802 38650
rect 13802 38598 13814 38650
rect 13814 38598 13844 38650
rect 13868 38598 13878 38650
rect 13878 38598 13924 38650
rect 13628 38596 13684 38598
rect 13708 38596 13764 38598
rect 13788 38596 13844 38598
rect 13868 38596 13924 38598
rect 9404 38106 9460 38108
rect 9484 38106 9540 38108
rect 9564 38106 9620 38108
rect 9644 38106 9700 38108
rect 9404 38054 9450 38106
rect 9450 38054 9460 38106
rect 9484 38054 9514 38106
rect 9514 38054 9526 38106
rect 9526 38054 9540 38106
rect 9564 38054 9578 38106
rect 9578 38054 9590 38106
rect 9590 38054 9620 38106
rect 9644 38054 9654 38106
rect 9654 38054 9700 38106
rect 9404 38052 9460 38054
rect 9484 38052 9540 38054
rect 9564 38052 9620 38054
rect 9644 38052 9700 38054
rect 9404 37018 9460 37020
rect 9484 37018 9540 37020
rect 9564 37018 9620 37020
rect 9644 37018 9700 37020
rect 9404 36966 9450 37018
rect 9450 36966 9460 37018
rect 9484 36966 9514 37018
rect 9514 36966 9526 37018
rect 9526 36966 9540 37018
rect 9564 36966 9578 37018
rect 9578 36966 9590 37018
rect 9590 36966 9620 37018
rect 9644 36966 9654 37018
rect 9654 36966 9700 37018
rect 9404 36964 9460 36966
rect 9484 36964 9540 36966
rect 9564 36964 9620 36966
rect 9644 36964 9700 36966
rect 9404 35930 9460 35932
rect 9484 35930 9540 35932
rect 9564 35930 9620 35932
rect 9644 35930 9700 35932
rect 9404 35878 9450 35930
rect 9450 35878 9460 35930
rect 9484 35878 9514 35930
rect 9514 35878 9526 35930
rect 9526 35878 9540 35930
rect 9564 35878 9578 35930
rect 9578 35878 9590 35930
rect 9590 35878 9620 35930
rect 9644 35878 9654 35930
rect 9654 35878 9700 35930
rect 9404 35876 9460 35878
rect 9484 35876 9540 35878
rect 9564 35876 9620 35878
rect 9644 35876 9700 35878
rect 9404 34842 9460 34844
rect 9484 34842 9540 34844
rect 9564 34842 9620 34844
rect 9644 34842 9700 34844
rect 9404 34790 9450 34842
rect 9450 34790 9460 34842
rect 9484 34790 9514 34842
rect 9514 34790 9526 34842
rect 9526 34790 9540 34842
rect 9564 34790 9578 34842
rect 9578 34790 9590 34842
rect 9590 34790 9620 34842
rect 9644 34790 9654 34842
rect 9654 34790 9700 34842
rect 9404 34788 9460 34790
rect 9484 34788 9540 34790
rect 9564 34788 9620 34790
rect 9644 34788 9700 34790
rect 9404 33754 9460 33756
rect 9484 33754 9540 33756
rect 9564 33754 9620 33756
rect 9644 33754 9700 33756
rect 9404 33702 9450 33754
rect 9450 33702 9460 33754
rect 9484 33702 9514 33754
rect 9514 33702 9526 33754
rect 9526 33702 9540 33754
rect 9564 33702 9578 33754
rect 9578 33702 9590 33754
rect 9590 33702 9620 33754
rect 9644 33702 9654 33754
rect 9654 33702 9700 33754
rect 9404 33700 9460 33702
rect 9484 33700 9540 33702
rect 9564 33700 9620 33702
rect 9644 33700 9700 33702
rect 9404 32666 9460 32668
rect 9484 32666 9540 32668
rect 9564 32666 9620 32668
rect 9644 32666 9700 32668
rect 9404 32614 9450 32666
rect 9450 32614 9460 32666
rect 9484 32614 9514 32666
rect 9514 32614 9526 32666
rect 9526 32614 9540 32666
rect 9564 32614 9578 32666
rect 9578 32614 9590 32666
rect 9590 32614 9620 32666
rect 9644 32614 9654 32666
rect 9654 32614 9700 32666
rect 9404 32612 9460 32614
rect 9484 32612 9540 32614
rect 9564 32612 9620 32614
rect 9644 32612 9700 32614
rect 9404 31578 9460 31580
rect 9484 31578 9540 31580
rect 9564 31578 9620 31580
rect 9644 31578 9700 31580
rect 9404 31526 9450 31578
rect 9450 31526 9460 31578
rect 9484 31526 9514 31578
rect 9514 31526 9526 31578
rect 9526 31526 9540 31578
rect 9564 31526 9578 31578
rect 9578 31526 9590 31578
rect 9590 31526 9620 31578
rect 9644 31526 9654 31578
rect 9654 31526 9700 31578
rect 9404 31524 9460 31526
rect 9484 31524 9540 31526
rect 9564 31524 9620 31526
rect 9644 31524 9700 31526
rect 9404 30490 9460 30492
rect 9484 30490 9540 30492
rect 9564 30490 9620 30492
rect 9644 30490 9700 30492
rect 9404 30438 9450 30490
rect 9450 30438 9460 30490
rect 9484 30438 9514 30490
rect 9514 30438 9526 30490
rect 9526 30438 9540 30490
rect 9564 30438 9578 30490
rect 9578 30438 9590 30490
rect 9590 30438 9620 30490
rect 9644 30438 9654 30490
rect 9654 30438 9700 30490
rect 9404 30436 9460 30438
rect 9484 30436 9540 30438
rect 9564 30436 9620 30438
rect 9644 30436 9700 30438
rect 9404 29402 9460 29404
rect 9484 29402 9540 29404
rect 9564 29402 9620 29404
rect 9644 29402 9700 29404
rect 9404 29350 9450 29402
rect 9450 29350 9460 29402
rect 9484 29350 9514 29402
rect 9514 29350 9526 29402
rect 9526 29350 9540 29402
rect 9564 29350 9578 29402
rect 9578 29350 9590 29402
rect 9590 29350 9620 29402
rect 9644 29350 9654 29402
rect 9654 29350 9700 29402
rect 9404 29348 9460 29350
rect 9484 29348 9540 29350
rect 9564 29348 9620 29350
rect 9644 29348 9700 29350
rect 9404 28314 9460 28316
rect 9484 28314 9540 28316
rect 9564 28314 9620 28316
rect 9644 28314 9700 28316
rect 9404 28262 9450 28314
rect 9450 28262 9460 28314
rect 9484 28262 9514 28314
rect 9514 28262 9526 28314
rect 9526 28262 9540 28314
rect 9564 28262 9578 28314
rect 9578 28262 9590 28314
rect 9590 28262 9620 28314
rect 9644 28262 9654 28314
rect 9654 28262 9700 28314
rect 9404 28260 9460 28262
rect 9484 28260 9540 28262
rect 9564 28260 9620 28262
rect 9644 28260 9700 28262
rect 9404 27226 9460 27228
rect 9484 27226 9540 27228
rect 9564 27226 9620 27228
rect 9644 27226 9700 27228
rect 9404 27174 9450 27226
rect 9450 27174 9460 27226
rect 9484 27174 9514 27226
rect 9514 27174 9526 27226
rect 9526 27174 9540 27226
rect 9564 27174 9578 27226
rect 9578 27174 9590 27226
rect 9590 27174 9620 27226
rect 9644 27174 9654 27226
rect 9654 27174 9700 27226
rect 9404 27172 9460 27174
rect 9484 27172 9540 27174
rect 9564 27172 9620 27174
rect 9644 27172 9700 27174
rect 9404 26138 9460 26140
rect 9484 26138 9540 26140
rect 9564 26138 9620 26140
rect 9644 26138 9700 26140
rect 9404 26086 9450 26138
rect 9450 26086 9460 26138
rect 9484 26086 9514 26138
rect 9514 26086 9526 26138
rect 9526 26086 9540 26138
rect 9564 26086 9578 26138
rect 9578 26086 9590 26138
rect 9590 26086 9620 26138
rect 9644 26086 9654 26138
rect 9654 26086 9700 26138
rect 9404 26084 9460 26086
rect 9484 26084 9540 26086
rect 9564 26084 9620 26086
rect 9644 26084 9700 26086
rect 4066 11600 4122 11656
rect 5180 12538 5236 12540
rect 5260 12538 5316 12540
rect 5340 12538 5396 12540
rect 5420 12538 5476 12540
rect 5180 12486 5226 12538
rect 5226 12486 5236 12538
rect 5260 12486 5290 12538
rect 5290 12486 5302 12538
rect 5302 12486 5316 12538
rect 5340 12486 5354 12538
rect 5354 12486 5366 12538
rect 5366 12486 5396 12538
rect 5420 12486 5430 12538
rect 5430 12486 5476 12538
rect 5180 12484 5236 12486
rect 5260 12484 5316 12486
rect 5340 12484 5396 12486
rect 5420 12484 5476 12486
rect 5180 11450 5236 11452
rect 5260 11450 5316 11452
rect 5340 11450 5396 11452
rect 5420 11450 5476 11452
rect 5180 11398 5226 11450
rect 5226 11398 5236 11450
rect 5260 11398 5290 11450
rect 5290 11398 5302 11450
rect 5302 11398 5316 11450
rect 5340 11398 5354 11450
rect 5354 11398 5366 11450
rect 5366 11398 5396 11450
rect 5420 11398 5430 11450
rect 5430 11398 5476 11450
rect 5180 11396 5236 11398
rect 5260 11396 5316 11398
rect 5340 11396 5396 11398
rect 5420 11396 5476 11398
rect 3146 8236 3148 8256
rect 3148 8236 3200 8256
rect 3200 8236 3202 8256
rect 3146 8200 3202 8236
rect 3146 7520 3202 7576
rect 2778 4800 2834 4856
rect 5180 10362 5236 10364
rect 5260 10362 5316 10364
rect 5340 10362 5396 10364
rect 5420 10362 5476 10364
rect 5180 10310 5226 10362
rect 5226 10310 5236 10362
rect 5260 10310 5290 10362
rect 5290 10310 5302 10362
rect 5302 10310 5316 10362
rect 5340 10310 5354 10362
rect 5354 10310 5366 10362
rect 5366 10310 5396 10362
rect 5420 10310 5430 10362
rect 5430 10310 5476 10362
rect 5180 10308 5236 10310
rect 5260 10308 5316 10310
rect 5340 10308 5396 10310
rect 5420 10308 5476 10310
rect 5180 9274 5236 9276
rect 5260 9274 5316 9276
rect 5340 9274 5396 9276
rect 5420 9274 5476 9276
rect 5180 9222 5226 9274
rect 5226 9222 5236 9274
rect 5260 9222 5290 9274
rect 5290 9222 5302 9274
rect 5302 9222 5316 9274
rect 5340 9222 5354 9274
rect 5354 9222 5366 9274
rect 5366 9222 5396 9274
rect 5420 9222 5430 9274
rect 5430 9222 5476 9274
rect 5180 9220 5236 9222
rect 5260 9220 5316 9222
rect 5340 9220 5396 9222
rect 5420 9220 5476 9222
rect 5180 8186 5236 8188
rect 5260 8186 5316 8188
rect 5340 8186 5396 8188
rect 5420 8186 5476 8188
rect 5180 8134 5226 8186
rect 5226 8134 5236 8186
rect 5260 8134 5290 8186
rect 5290 8134 5302 8186
rect 5302 8134 5316 8186
rect 5340 8134 5354 8186
rect 5354 8134 5366 8186
rect 5366 8134 5396 8186
rect 5420 8134 5430 8186
rect 5430 8134 5476 8186
rect 5180 8132 5236 8134
rect 5260 8132 5316 8134
rect 5340 8132 5396 8134
rect 5420 8132 5476 8134
rect 5180 7098 5236 7100
rect 5260 7098 5316 7100
rect 5340 7098 5396 7100
rect 5420 7098 5476 7100
rect 5180 7046 5226 7098
rect 5226 7046 5236 7098
rect 5260 7046 5290 7098
rect 5290 7046 5302 7098
rect 5302 7046 5316 7098
rect 5340 7046 5354 7098
rect 5354 7046 5366 7098
rect 5366 7046 5396 7098
rect 5420 7046 5430 7098
rect 5430 7046 5476 7098
rect 5180 7044 5236 7046
rect 5260 7044 5316 7046
rect 5340 7044 5396 7046
rect 5420 7044 5476 7046
rect 5180 6010 5236 6012
rect 5260 6010 5316 6012
rect 5340 6010 5396 6012
rect 5420 6010 5476 6012
rect 5180 5958 5226 6010
rect 5226 5958 5236 6010
rect 5260 5958 5290 6010
rect 5290 5958 5302 6010
rect 5302 5958 5316 6010
rect 5340 5958 5354 6010
rect 5354 5958 5366 6010
rect 5366 5958 5396 6010
rect 5420 5958 5430 6010
rect 5430 5958 5476 6010
rect 5180 5956 5236 5958
rect 5260 5956 5316 5958
rect 5340 5956 5396 5958
rect 5420 5956 5476 5958
rect 3422 5480 3478 5536
rect 5180 4922 5236 4924
rect 5260 4922 5316 4924
rect 5340 4922 5396 4924
rect 5420 4922 5476 4924
rect 5180 4870 5226 4922
rect 5226 4870 5236 4922
rect 5260 4870 5290 4922
rect 5290 4870 5302 4922
rect 5302 4870 5316 4922
rect 5340 4870 5354 4922
rect 5354 4870 5366 4922
rect 5366 4870 5396 4922
rect 5420 4870 5430 4922
rect 5430 4870 5476 4922
rect 5180 4868 5236 4870
rect 5260 4868 5316 4870
rect 5340 4868 5396 4870
rect 5420 4868 5476 4870
rect 3422 4120 3478 4176
rect 3422 3440 3478 3496
rect 3422 2760 3478 2816
rect 3422 2080 3478 2136
rect 3330 1400 3386 1456
rect 5180 3834 5236 3836
rect 5260 3834 5316 3836
rect 5340 3834 5396 3836
rect 5420 3834 5476 3836
rect 5180 3782 5226 3834
rect 5226 3782 5236 3834
rect 5260 3782 5290 3834
rect 5290 3782 5302 3834
rect 5302 3782 5316 3834
rect 5340 3782 5354 3834
rect 5354 3782 5366 3834
rect 5366 3782 5396 3834
rect 5420 3782 5430 3834
rect 5430 3782 5476 3834
rect 5180 3780 5236 3782
rect 5260 3780 5316 3782
rect 5340 3780 5396 3782
rect 5420 3780 5476 3782
rect 5180 2746 5236 2748
rect 5260 2746 5316 2748
rect 5340 2746 5396 2748
rect 5420 2746 5476 2748
rect 5180 2694 5226 2746
rect 5226 2694 5236 2746
rect 5260 2694 5290 2746
rect 5290 2694 5302 2746
rect 5302 2694 5316 2746
rect 5340 2694 5354 2746
rect 5354 2694 5366 2746
rect 5366 2694 5396 2746
rect 5420 2694 5430 2746
rect 5430 2694 5476 2746
rect 5180 2692 5236 2694
rect 5260 2692 5316 2694
rect 5340 2692 5396 2694
rect 5420 2692 5476 2694
rect 9404 25050 9460 25052
rect 9484 25050 9540 25052
rect 9564 25050 9620 25052
rect 9644 25050 9700 25052
rect 9404 24998 9450 25050
rect 9450 24998 9460 25050
rect 9484 24998 9514 25050
rect 9514 24998 9526 25050
rect 9526 24998 9540 25050
rect 9564 24998 9578 25050
rect 9578 24998 9590 25050
rect 9590 24998 9620 25050
rect 9644 24998 9654 25050
rect 9654 24998 9700 25050
rect 9404 24996 9460 24998
rect 9484 24996 9540 24998
rect 9564 24996 9620 24998
rect 9644 24996 9700 24998
rect 9404 23962 9460 23964
rect 9484 23962 9540 23964
rect 9564 23962 9620 23964
rect 9644 23962 9700 23964
rect 9404 23910 9450 23962
rect 9450 23910 9460 23962
rect 9484 23910 9514 23962
rect 9514 23910 9526 23962
rect 9526 23910 9540 23962
rect 9564 23910 9578 23962
rect 9578 23910 9590 23962
rect 9590 23910 9620 23962
rect 9644 23910 9654 23962
rect 9654 23910 9700 23962
rect 9404 23908 9460 23910
rect 9484 23908 9540 23910
rect 9564 23908 9620 23910
rect 9644 23908 9700 23910
rect 9404 22874 9460 22876
rect 9484 22874 9540 22876
rect 9564 22874 9620 22876
rect 9644 22874 9700 22876
rect 9404 22822 9450 22874
rect 9450 22822 9460 22874
rect 9484 22822 9514 22874
rect 9514 22822 9526 22874
rect 9526 22822 9540 22874
rect 9564 22822 9578 22874
rect 9578 22822 9590 22874
rect 9590 22822 9620 22874
rect 9644 22822 9654 22874
rect 9654 22822 9700 22874
rect 9404 22820 9460 22822
rect 9484 22820 9540 22822
rect 9564 22820 9620 22822
rect 9644 22820 9700 22822
rect 9404 21786 9460 21788
rect 9484 21786 9540 21788
rect 9564 21786 9620 21788
rect 9644 21786 9700 21788
rect 9404 21734 9450 21786
rect 9450 21734 9460 21786
rect 9484 21734 9514 21786
rect 9514 21734 9526 21786
rect 9526 21734 9540 21786
rect 9564 21734 9578 21786
rect 9578 21734 9590 21786
rect 9590 21734 9620 21786
rect 9644 21734 9654 21786
rect 9654 21734 9700 21786
rect 9404 21732 9460 21734
rect 9484 21732 9540 21734
rect 9564 21732 9620 21734
rect 9644 21732 9700 21734
rect 9404 20698 9460 20700
rect 9484 20698 9540 20700
rect 9564 20698 9620 20700
rect 9644 20698 9700 20700
rect 9404 20646 9450 20698
rect 9450 20646 9460 20698
rect 9484 20646 9514 20698
rect 9514 20646 9526 20698
rect 9526 20646 9540 20698
rect 9564 20646 9578 20698
rect 9578 20646 9590 20698
rect 9590 20646 9620 20698
rect 9644 20646 9654 20698
rect 9654 20646 9700 20698
rect 9404 20644 9460 20646
rect 9484 20644 9540 20646
rect 9564 20644 9620 20646
rect 9644 20644 9700 20646
rect 13628 37562 13684 37564
rect 13708 37562 13764 37564
rect 13788 37562 13844 37564
rect 13868 37562 13924 37564
rect 13628 37510 13674 37562
rect 13674 37510 13684 37562
rect 13708 37510 13738 37562
rect 13738 37510 13750 37562
rect 13750 37510 13764 37562
rect 13788 37510 13802 37562
rect 13802 37510 13814 37562
rect 13814 37510 13844 37562
rect 13868 37510 13878 37562
rect 13878 37510 13924 37562
rect 13628 37508 13684 37510
rect 13708 37508 13764 37510
rect 13788 37508 13844 37510
rect 13868 37508 13924 37510
rect 13628 36474 13684 36476
rect 13708 36474 13764 36476
rect 13788 36474 13844 36476
rect 13868 36474 13924 36476
rect 13628 36422 13674 36474
rect 13674 36422 13684 36474
rect 13708 36422 13738 36474
rect 13738 36422 13750 36474
rect 13750 36422 13764 36474
rect 13788 36422 13802 36474
rect 13802 36422 13814 36474
rect 13814 36422 13844 36474
rect 13868 36422 13878 36474
rect 13878 36422 13924 36474
rect 13628 36420 13684 36422
rect 13708 36420 13764 36422
rect 13788 36420 13844 36422
rect 13868 36420 13924 36422
rect 13628 35386 13684 35388
rect 13708 35386 13764 35388
rect 13788 35386 13844 35388
rect 13868 35386 13924 35388
rect 13628 35334 13674 35386
rect 13674 35334 13684 35386
rect 13708 35334 13738 35386
rect 13738 35334 13750 35386
rect 13750 35334 13764 35386
rect 13788 35334 13802 35386
rect 13802 35334 13814 35386
rect 13814 35334 13844 35386
rect 13868 35334 13878 35386
rect 13878 35334 13924 35386
rect 13628 35332 13684 35334
rect 13708 35332 13764 35334
rect 13788 35332 13844 35334
rect 13868 35332 13924 35334
rect 13628 34298 13684 34300
rect 13708 34298 13764 34300
rect 13788 34298 13844 34300
rect 13868 34298 13924 34300
rect 13628 34246 13674 34298
rect 13674 34246 13684 34298
rect 13708 34246 13738 34298
rect 13738 34246 13750 34298
rect 13750 34246 13764 34298
rect 13788 34246 13802 34298
rect 13802 34246 13814 34298
rect 13814 34246 13844 34298
rect 13868 34246 13878 34298
rect 13878 34246 13924 34298
rect 13628 34244 13684 34246
rect 13708 34244 13764 34246
rect 13788 34244 13844 34246
rect 13868 34244 13924 34246
rect 13628 33210 13684 33212
rect 13708 33210 13764 33212
rect 13788 33210 13844 33212
rect 13868 33210 13924 33212
rect 13628 33158 13674 33210
rect 13674 33158 13684 33210
rect 13708 33158 13738 33210
rect 13738 33158 13750 33210
rect 13750 33158 13764 33210
rect 13788 33158 13802 33210
rect 13802 33158 13814 33210
rect 13814 33158 13844 33210
rect 13868 33158 13878 33210
rect 13878 33158 13924 33210
rect 13628 33156 13684 33158
rect 13708 33156 13764 33158
rect 13788 33156 13844 33158
rect 13868 33156 13924 33158
rect 13628 32122 13684 32124
rect 13708 32122 13764 32124
rect 13788 32122 13844 32124
rect 13868 32122 13924 32124
rect 13628 32070 13674 32122
rect 13674 32070 13684 32122
rect 13708 32070 13738 32122
rect 13738 32070 13750 32122
rect 13750 32070 13764 32122
rect 13788 32070 13802 32122
rect 13802 32070 13814 32122
rect 13814 32070 13844 32122
rect 13868 32070 13878 32122
rect 13878 32070 13924 32122
rect 13628 32068 13684 32070
rect 13708 32068 13764 32070
rect 13788 32068 13844 32070
rect 13868 32068 13924 32070
rect 13628 31034 13684 31036
rect 13708 31034 13764 31036
rect 13788 31034 13844 31036
rect 13868 31034 13924 31036
rect 13628 30982 13674 31034
rect 13674 30982 13684 31034
rect 13708 30982 13738 31034
rect 13738 30982 13750 31034
rect 13750 30982 13764 31034
rect 13788 30982 13802 31034
rect 13802 30982 13814 31034
rect 13814 30982 13844 31034
rect 13868 30982 13878 31034
rect 13878 30982 13924 31034
rect 13628 30980 13684 30982
rect 13708 30980 13764 30982
rect 13788 30980 13844 30982
rect 13868 30980 13924 30982
rect 17852 39194 17908 39196
rect 17932 39194 17988 39196
rect 18012 39194 18068 39196
rect 18092 39194 18148 39196
rect 17852 39142 17898 39194
rect 17898 39142 17908 39194
rect 17932 39142 17962 39194
rect 17962 39142 17974 39194
rect 17974 39142 17988 39194
rect 18012 39142 18026 39194
rect 18026 39142 18038 39194
rect 18038 39142 18068 39194
rect 18092 39142 18102 39194
rect 18102 39142 18148 39194
rect 17852 39140 17908 39142
rect 17932 39140 17988 39142
rect 18012 39140 18068 39142
rect 18092 39140 18148 39142
rect 17852 38106 17908 38108
rect 17932 38106 17988 38108
rect 18012 38106 18068 38108
rect 18092 38106 18148 38108
rect 17852 38054 17898 38106
rect 17898 38054 17908 38106
rect 17932 38054 17962 38106
rect 17962 38054 17974 38106
rect 17974 38054 17988 38106
rect 18012 38054 18026 38106
rect 18026 38054 18038 38106
rect 18038 38054 18068 38106
rect 18092 38054 18102 38106
rect 18102 38054 18148 38106
rect 17852 38052 17908 38054
rect 17932 38052 17988 38054
rect 18012 38052 18068 38054
rect 18092 38052 18148 38054
rect 17852 37018 17908 37020
rect 17932 37018 17988 37020
rect 18012 37018 18068 37020
rect 18092 37018 18148 37020
rect 17852 36966 17898 37018
rect 17898 36966 17908 37018
rect 17932 36966 17962 37018
rect 17962 36966 17974 37018
rect 17974 36966 17988 37018
rect 18012 36966 18026 37018
rect 18026 36966 18038 37018
rect 18038 36966 18068 37018
rect 18092 36966 18102 37018
rect 18102 36966 18148 37018
rect 17852 36964 17908 36966
rect 17932 36964 17988 36966
rect 18012 36964 18068 36966
rect 18092 36964 18148 36966
rect 13628 29946 13684 29948
rect 13708 29946 13764 29948
rect 13788 29946 13844 29948
rect 13868 29946 13924 29948
rect 13628 29894 13674 29946
rect 13674 29894 13684 29946
rect 13708 29894 13738 29946
rect 13738 29894 13750 29946
rect 13750 29894 13764 29946
rect 13788 29894 13802 29946
rect 13802 29894 13814 29946
rect 13814 29894 13844 29946
rect 13868 29894 13878 29946
rect 13878 29894 13924 29946
rect 13628 29892 13684 29894
rect 13708 29892 13764 29894
rect 13788 29892 13844 29894
rect 13868 29892 13924 29894
rect 13628 28858 13684 28860
rect 13708 28858 13764 28860
rect 13788 28858 13844 28860
rect 13868 28858 13924 28860
rect 13628 28806 13674 28858
rect 13674 28806 13684 28858
rect 13708 28806 13738 28858
rect 13738 28806 13750 28858
rect 13750 28806 13764 28858
rect 13788 28806 13802 28858
rect 13802 28806 13814 28858
rect 13814 28806 13844 28858
rect 13868 28806 13878 28858
rect 13878 28806 13924 28858
rect 13628 28804 13684 28806
rect 13708 28804 13764 28806
rect 13788 28804 13844 28806
rect 13868 28804 13924 28806
rect 13628 27770 13684 27772
rect 13708 27770 13764 27772
rect 13788 27770 13844 27772
rect 13868 27770 13924 27772
rect 13628 27718 13674 27770
rect 13674 27718 13684 27770
rect 13708 27718 13738 27770
rect 13738 27718 13750 27770
rect 13750 27718 13764 27770
rect 13788 27718 13802 27770
rect 13802 27718 13814 27770
rect 13814 27718 13844 27770
rect 13868 27718 13878 27770
rect 13878 27718 13924 27770
rect 13628 27716 13684 27718
rect 13708 27716 13764 27718
rect 13788 27716 13844 27718
rect 13868 27716 13924 27718
rect 13628 26682 13684 26684
rect 13708 26682 13764 26684
rect 13788 26682 13844 26684
rect 13868 26682 13924 26684
rect 13628 26630 13674 26682
rect 13674 26630 13684 26682
rect 13708 26630 13738 26682
rect 13738 26630 13750 26682
rect 13750 26630 13764 26682
rect 13788 26630 13802 26682
rect 13802 26630 13814 26682
rect 13814 26630 13844 26682
rect 13868 26630 13878 26682
rect 13878 26630 13924 26682
rect 13628 26628 13684 26630
rect 13708 26628 13764 26630
rect 13788 26628 13844 26630
rect 13868 26628 13924 26630
rect 13628 25594 13684 25596
rect 13708 25594 13764 25596
rect 13788 25594 13844 25596
rect 13868 25594 13924 25596
rect 13628 25542 13674 25594
rect 13674 25542 13684 25594
rect 13708 25542 13738 25594
rect 13738 25542 13750 25594
rect 13750 25542 13764 25594
rect 13788 25542 13802 25594
rect 13802 25542 13814 25594
rect 13814 25542 13844 25594
rect 13868 25542 13878 25594
rect 13878 25542 13924 25594
rect 13628 25540 13684 25542
rect 13708 25540 13764 25542
rect 13788 25540 13844 25542
rect 13868 25540 13924 25542
rect 13628 24506 13684 24508
rect 13708 24506 13764 24508
rect 13788 24506 13844 24508
rect 13868 24506 13924 24508
rect 13628 24454 13674 24506
rect 13674 24454 13684 24506
rect 13708 24454 13738 24506
rect 13738 24454 13750 24506
rect 13750 24454 13764 24506
rect 13788 24454 13802 24506
rect 13802 24454 13814 24506
rect 13814 24454 13844 24506
rect 13868 24454 13878 24506
rect 13878 24454 13924 24506
rect 13628 24452 13684 24454
rect 13708 24452 13764 24454
rect 13788 24452 13844 24454
rect 13868 24452 13924 24454
rect 9404 19610 9460 19612
rect 9484 19610 9540 19612
rect 9564 19610 9620 19612
rect 9644 19610 9700 19612
rect 9404 19558 9450 19610
rect 9450 19558 9460 19610
rect 9484 19558 9514 19610
rect 9514 19558 9526 19610
rect 9526 19558 9540 19610
rect 9564 19558 9578 19610
rect 9578 19558 9590 19610
rect 9590 19558 9620 19610
rect 9644 19558 9654 19610
rect 9654 19558 9700 19610
rect 9404 19556 9460 19558
rect 9484 19556 9540 19558
rect 9564 19556 9620 19558
rect 9644 19556 9700 19558
rect 9404 18522 9460 18524
rect 9484 18522 9540 18524
rect 9564 18522 9620 18524
rect 9644 18522 9700 18524
rect 9404 18470 9450 18522
rect 9450 18470 9460 18522
rect 9484 18470 9514 18522
rect 9514 18470 9526 18522
rect 9526 18470 9540 18522
rect 9564 18470 9578 18522
rect 9578 18470 9590 18522
rect 9590 18470 9620 18522
rect 9644 18470 9654 18522
rect 9654 18470 9700 18522
rect 9404 18468 9460 18470
rect 9484 18468 9540 18470
rect 9564 18468 9620 18470
rect 9644 18468 9700 18470
rect 9404 17434 9460 17436
rect 9484 17434 9540 17436
rect 9564 17434 9620 17436
rect 9644 17434 9700 17436
rect 9404 17382 9450 17434
rect 9450 17382 9460 17434
rect 9484 17382 9514 17434
rect 9514 17382 9526 17434
rect 9526 17382 9540 17434
rect 9564 17382 9578 17434
rect 9578 17382 9590 17434
rect 9590 17382 9620 17434
rect 9644 17382 9654 17434
rect 9654 17382 9700 17434
rect 9404 17380 9460 17382
rect 9484 17380 9540 17382
rect 9564 17380 9620 17382
rect 9644 17380 9700 17382
rect 9404 16346 9460 16348
rect 9484 16346 9540 16348
rect 9564 16346 9620 16348
rect 9644 16346 9700 16348
rect 9404 16294 9450 16346
rect 9450 16294 9460 16346
rect 9484 16294 9514 16346
rect 9514 16294 9526 16346
rect 9526 16294 9540 16346
rect 9564 16294 9578 16346
rect 9578 16294 9590 16346
rect 9590 16294 9620 16346
rect 9644 16294 9654 16346
rect 9654 16294 9700 16346
rect 9404 16292 9460 16294
rect 9484 16292 9540 16294
rect 9564 16292 9620 16294
rect 9644 16292 9700 16294
rect 9404 15258 9460 15260
rect 9484 15258 9540 15260
rect 9564 15258 9620 15260
rect 9644 15258 9700 15260
rect 9404 15206 9450 15258
rect 9450 15206 9460 15258
rect 9484 15206 9514 15258
rect 9514 15206 9526 15258
rect 9526 15206 9540 15258
rect 9564 15206 9578 15258
rect 9578 15206 9590 15258
rect 9590 15206 9620 15258
rect 9644 15206 9654 15258
rect 9654 15206 9700 15258
rect 9404 15204 9460 15206
rect 9484 15204 9540 15206
rect 9564 15204 9620 15206
rect 9644 15204 9700 15206
rect 9404 14170 9460 14172
rect 9484 14170 9540 14172
rect 9564 14170 9620 14172
rect 9644 14170 9700 14172
rect 9404 14118 9450 14170
rect 9450 14118 9460 14170
rect 9484 14118 9514 14170
rect 9514 14118 9526 14170
rect 9526 14118 9540 14170
rect 9564 14118 9578 14170
rect 9578 14118 9590 14170
rect 9590 14118 9620 14170
rect 9644 14118 9654 14170
rect 9654 14118 9700 14170
rect 9404 14116 9460 14118
rect 9484 14116 9540 14118
rect 9564 14116 9620 14118
rect 9644 14116 9700 14118
rect 9404 13082 9460 13084
rect 9484 13082 9540 13084
rect 9564 13082 9620 13084
rect 9644 13082 9700 13084
rect 9404 13030 9450 13082
rect 9450 13030 9460 13082
rect 9484 13030 9514 13082
rect 9514 13030 9526 13082
rect 9526 13030 9540 13082
rect 9564 13030 9578 13082
rect 9578 13030 9590 13082
rect 9590 13030 9620 13082
rect 9644 13030 9654 13082
rect 9654 13030 9700 13082
rect 9404 13028 9460 13030
rect 9484 13028 9540 13030
rect 9564 13028 9620 13030
rect 9644 13028 9700 13030
rect 9404 11994 9460 11996
rect 9484 11994 9540 11996
rect 9564 11994 9620 11996
rect 9644 11994 9700 11996
rect 9404 11942 9450 11994
rect 9450 11942 9460 11994
rect 9484 11942 9514 11994
rect 9514 11942 9526 11994
rect 9526 11942 9540 11994
rect 9564 11942 9578 11994
rect 9578 11942 9590 11994
rect 9590 11942 9620 11994
rect 9644 11942 9654 11994
rect 9654 11942 9700 11994
rect 9404 11940 9460 11942
rect 9484 11940 9540 11942
rect 9564 11940 9620 11942
rect 9644 11940 9700 11942
rect 9404 10906 9460 10908
rect 9484 10906 9540 10908
rect 9564 10906 9620 10908
rect 9644 10906 9700 10908
rect 9404 10854 9450 10906
rect 9450 10854 9460 10906
rect 9484 10854 9514 10906
rect 9514 10854 9526 10906
rect 9526 10854 9540 10906
rect 9564 10854 9578 10906
rect 9578 10854 9590 10906
rect 9590 10854 9620 10906
rect 9644 10854 9654 10906
rect 9654 10854 9700 10906
rect 9404 10852 9460 10854
rect 9484 10852 9540 10854
rect 9564 10852 9620 10854
rect 9644 10852 9700 10854
rect 9404 9818 9460 9820
rect 9484 9818 9540 9820
rect 9564 9818 9620 9820
rect 9644 9818 9700 9820
rect 9404 9766 9450 9818
rect 9450 9766 9460 9818
rect 9484 9766 9514 9818
rect 9514 9766 9526 9818
rect 9526 9766 9540 9818
rect 9564 9766 9578 9818
rect 9578 9766 9590 9818
rect 9590 9766 9620 9818
rect 9644 9766 9654 9818
rect 9654 9766 9700 9818
rect 9404 9764 9460 9766
rect 9484 9764 9540 9766
rect 9564 9764 9620 9766
rect 9644 9764 9700 9766
rect 9404 8730 9460 8732
rect 9484 8730 9540 8732
rect 9564 8730 9620 8732
rect 9644 8730 9700 8732
rect 9404 8678 9450 8730
rect 9450 8678 9460 8730
rect 9484 8678 9514 8730
rect 9514 8678 9526 8730
rect 9526 8678 9540 8730
rect 9564 8678 9578 8730
rect 9578 8678 9590 8730
rect 9590 8678 9620 8730
rect 9644 8678 9654 8730
rect 9654 8678 9700 8730
rect 9404 8676 9460 8678
rect 9484 8676 9540 8678
rect 9564 8676 9620 8678
rect 9644 8676 9700 8678
rect 9404 7642 9460 7644
rect 9484 7642 9540 7644
rect 9564 7642 9620 7644
rect 9644 7642 9700 7644
rect 9404 7590 9450 7642
rect 9450 7590 9460 7642
rect 9484 7590 9514 7642
rect 9514 7590 9526 7642
rect 9526 7590 9540 7642
rect 9564 7590 9578 7642
rect 9578 7590 9590 7642
rect 9590 7590 9620 7642
rect 9644 7590 9654 7642
rect 9654 7590 9700 7642
rect 9404 7588 9460 7590
rect 9484 7588 9540 7590
rect 9564 7588 9620 7590
rect 9644 7588 9700 7590
rect 9404 6554 9460 6556
rect 9484 6554 9540 6556
rect 9564 6554 9620 6556
rect 9644 6554 9700 6556
rect 9404 6502 9450 6554
rect 9450 6502 9460 6554
rect 9484 6502 9514 6554
rect 9514 6502 9526 6554
rect 9526 6502 9540 6554
rect 9564 6502 9578 6554
rect 9578 6502 9590 6554
rect 9590 6502 9620 6554
rect 9644 6502 9654 6554
rect 9654 6502 9700 6554
rect 9404 6500 9460 6502
rect 9484 6500 9540 6502
rect 9564 6500 9620 6502
rect 9644 6500 9700 6502
rect 9404 5466 9460 5468
rect 9484 5466 9540 5468
rect 9564 5466 9620 5468
rect 9644 5466 9700 5468
rect 9404 5414 9450 5466
rect 9450 5414 9460 5466
rect 9484 5414 9514 5466
rect 9514 5414 9526 5466
rect 9526 5414 9540 5466
rect 9564 5414 9578 5466
rect 9578 5414 9590 5466
rect 9590 5414 9620 5466
rect 9644 5414 9654 5466
rect 9654 5414 9700 5466
rect 9404 5412 9460 5414
rect 9484 5412 9540 5414
rect 9564 5412 9620 5414
rect 9644 5412 9700 5414
rect 9404 4378 9460 4380
rect 9484 4378 9540 4380
rect 9564 4378 9620 4380
rect 9644 4378 9700 4380
rect 9404 4326 9450 4378
rect 9450 4326 9460 4378
rect 9484 4326 9514 4378
rect 9514 4326 9526 4378
rect 9526 4326 9540 4378
rect 9564 4326 9578 4378
rect 9578 4326 9590 4378
rect 9590 4326 9620 4378
rect 9644 4326 9654 4378
rect 9654 4326 9700 4378
rect 9404 4324 9460 4326
rect 9484 4324 9540 4326
rect 9564 4324 9620 4326
rect 9644 4324 9700 4326
rect 9404 3290 9460 3292
rect 9484 3290 9540 3292
rect 9564 3290 9620 3292
rect 9644 3290 9700 3292
rect 9404 3238 9450 3290
rect 9450 3238 9460 3290
rect 9484 3238 9514 3290
rect 9514 3238 9526 3290
rect 9526 3238 9540 3290
rect 9564 3238 9578 3290
rect 9578 3238 9590 3290
rect 9590 3238 9620 3290
rect 9644 3238 9654 3290
rect 9654 3238 9700 3290
rect 9404 3236 9460 3238
rect 9484 3236 9540 3238
rect 9564 3236 9620 3238
rect 9644 3236 9700 3238
rect 9404 2202 9460 2204
rect 9484 2202 9540 2204
rect 9564 2202 9620 2204
rect 9644 2202 9700 2204
rect 9404 2150 9450 2202
rect 9450 2150 9460 2202
rect 9484 2150 9514 2202
rect 9514 2150 9526 2202
rect 9526 2150 9540 2202
rect 9564 2150 9578 2202
rect 9578 2150 9590 2202
rect 9590 2150 9620 2202
rect 9644 2150 9654 2202
rect 9654 2150 9700 2202
rect 9404 2148 9460 2150
rect 9484 2148 9540 2150
rect 9564 2148 9620 2150
rect 9644 2148 9700 2150
rect 13628 23418 13684 23420
rect 13708 23418 13764 23420
rect 13788 23418 13844 23420
rect 13868 23418 13924 23420
rect 13628 23366 13674 23418
rect 13674 23366 13684 23418
rect 13708 23366 13738 23418
rect 13738 23366 13750 23418
rect 13750 23366 13764 23418
rect 13788 23366 13802 23418
rect 13802 23366 13814 23418
rect 13814 23366 13844 23418
rect 13868 23366 13878 23418
rect 13878 23366 13924 23418
rect 13628 23364 13684 23366
rect 13708 23364 13764 23366
rect 13788 23364 13844 23366
rect 13868 23364 13924 23366
rect 13628 22330 13684 22332
rect 13708 22330 13764 22332
rect 13788 22330 13844 22332
rect 13868 22330 13924 22332
rect 13628 22278 13674 22330
rect 13674 22278 13684 22330
rect 13708 22278 13738 22330
rect 13738 22278 13750 22330
rect 13750 22278 13764 22330
rect 13788 22278 13802 22330
rect 13802 22278 13814 22330
rect 13814 22278 13844 22330
rect 13868 22278 13878 22330
rect 13878 22278 13924 22330
rect 13628 22276 13684 22278
rect 13708 22276 13764 22278
rect 13788 22276 13844 22278
rect 13868 22276 13924 22278
rect 13628 21242 13684 21244
rect 13708 21242 13764 21244
rect 13788 21242 13844 21244
rect 13868 21242 13924 21244
rect 13628 21190 13674 21242
rect 13674 21190 13684 21242
rect 13708 21190 13738 21242
rect 13738 21190 13750 21242
rect 13750 21190 13764 21242
rect 13788 21190 13802 21242
rect 13802 21190 13814 21242
rect 13814 21190 13844 21242
rect 13868 21190 13878 21242
rect 13878 21190 13924 21242
rect 13628 21188 13684 21190
rect 13708 21188 13764 21190
rect 13788 21188 13844 21190
rect 13868 21188 13924 21190
rect 13628 20154 13684 20156
rect 13708 20154 13764 20156
rect 13788 20154 13844 20156
rect 13868 20154 13924 20156
rect 13628 20102 13674 20154
rect 13674 20102 13684 20154
rect 13708 20102 13738 20154
rect 13738 20102 13750 20154
rect 13750 20102 13764 20154
rect 13788 20102 13802 20154
rect 13802 20102 13814 20154
rect 13814 20102 13844 20154
rect 13868 20102 13878 20154
rect 13878 20102 13924 20154
rect 13628 20100 13684 20102
rect 13708 20100 13764 20102
rect 13788 20100 13844 20102
rect 13868 20100 13924 20102
rect 17852 35930 17908 35932
rect 17932 35930 17988 35932
rect 18012 35930 18068 35932
rect 18092 35930 18148 35932
rect 17852 35878 17898 35930
rect 17898 35878 17908 35930
rect 17932 35878 17962 35930
rect 17962 35878 17974 35930
rect 17974 35878 17988 35930
rect 18012 35878 18026 35930
rect 18026 35878 18038 35930
rect 18038 35878 18068 35930
rect 18092 35878 18102 35930
rect 18102 35878 18148 35930
rect 17852 35876 17908 35878
rect 17932 35876 17988 35878
rect 18012 35876 18068 35878
rect 18092 35876 18148 35878
rect 22076 39738 22132 39740
rect 22156 39738 22212 39740
rect 22236 39738 22292 39740
rect 22316 39738 22372 39740
rect 22076 39686 22122 39738
rect 22122 39686 22132 39738
rect 22156 39686 22186 39738
rect 22186 39686 22198 39738
rect 22198 39686 22212 39738
rect 22236 39686 22250 39738
rect 22250 39686 22262 39738
rect 22262 39686 22292 39738
rect 22316 39686 22326 39738
rect 22326 39686 22372 39738
rect 22076 39684 22132 39686
rect 22156 39684 22212 39686
rect 22236 39684 22292 39686
rect 22316 39684 22372 39686
rect 17852 34842 17908 34844
rect 17932 34842 17988 34844
rect 18012 34842 18068 34844
rect 18092 34842 18148 34844
rect 17852 34790 17898 34842
rect 17898 34790 17908 34842
rect 17932 34790 17962 34842
rect 17962 34790 17974 34842
rect 17974 34790 17988 34842
rect 18012 34790 18026 34842
rect 18026 34790 18038 34842
rect 18038 34790 18068 34842
rect 18092 34790 18102 34842
rect 18102 34790 18148 34842
rect 17852 34788 17908 34790
rect 17932 34788 17988 34790
rect 18012 34788 18068 34790
rect 18092 34788 18148 34790
rect 17852 33754 17908 33756
rect 17932 33754 17988 33756
rect 18012 33754 18068 33756
rect 18092 33754 18148 33756
rect 17852 33702 17898 33754
rect 17898 33702 17908 33754
rect 17932 33702 17962 33754
rect 17962 33702 17974 33754
rect 17974 33702 17988 33754
rect 18012 33702 18026 33754
rect 18026 33702 18038 33754
rect 18038 33702 18068 33754
rect 18092 33702 18102 33754
rect 18102 33702 18148 33754
rect 17852 33700 17908 33702
rect 17932 33700 17988 33702
rect 18012 33700 18068 33702
rect 18092 33700 18148 33702
rect 17852 32666 17908 32668
rect 17932 32666 17988 32668
rect 18012 32666 18068 32668
rect 18092 32666 18148 32668
rect 17852 32614 17898 32666
rect 17898 32614 17908 32666
rect 17932 32614 17962 32666
rect 17962 32614 17974 32666
rect 17974 32614 17988 32666
rect 18012 32614 18026 32666
rect 18026 32614 18038 32666
rect 18038 32614 18068 32666
rect 18092 32614 18102 32666
rect 18102 32614 18148 32666
rect 17852 32612 17908 32614
rect 17932 32612 17988 32614
rect 18012 32612 18068 32614
rect 18092 32612 18148 32614
rect 22076 38650 22132 38652
rect 22156 38650 22212 38652
rect 22236 38650 22292 38652
rect 22316 38650 22372 38652
rect 22076 38598 22122 38650
rect 22122 38598 22132 38650
rect 22156 38598 22186 38650
rect 22186 38598 22198 38650
rect 22198 38598 22212 38650
rect 22236 38598 22250 38650
rect 22250 38598 22262 38650
rect 22262 38598 22292 38650
rect 22316 38598 22326 38650
rect 22326 38598 22372 38650
rect 22076 38596 22132 38598
rect 22156 38596 22212 38598
rect 22236 38596 22292 38598
rect 22316 38596 22372 38598
rect 22076 37562 22132 37564
rect 22156 37562 22212 37564
rect 22236 37562 22292 37564
rect 22316 37562 22372 37564
rect 22076 37510 22122 37562
rect 22122 37510 22132 37562
rect 22156 37510 22186 37562
rect 22186 37510 22198 37562
rect 22198 37510 22212 37562
rect 22236 37510 22250 37562
rect 22250 37510 22262 37562
rect 22262 37510 22292 37562
rect 22316 37510 22326 37562
rect 22326 37510 22372 37562
rect 22076 37508 22132 37510
rect 22156 37508 22212 37510
rect 22236 37508 22292 37510
rect 22316 37508 22372 37510
rect 22076 36474 22132 36476
rect 22156 36474 22212 36476
rect 22236 36474 22292 36476
rect 22316 36474 22372 36476
rect 22076 36422 22122 36474
rect 22122 36422 22132 36474
rect 22156 36422 22186 36474
rect 22186 36422 22198 36474
rect 22198 36422 22212 36474
rect 22236 36422 22250 36474
rect 22250 36422 22262 36474
rect 22262 36422 22292 36474
rect 22316 36422 22326 36474
rect 22326 36422 22372 36474
rect 22076 36420 22132 36422
rect 22156 36420 22212 36422
rect 22236 36420 22292 36422
rect 22316 36420 22372 36422
rect 22076 35386 22132 35388
rect 22156 35386 22212 35388
rect 22236 35386 22292 35388
rect 22316 35386 22372 35388
rect 22076 35334 22122 35386
rect 22122 35334 22132 35386
rect 22156 35334 22186 35386
rect 22186 35334 22198 35386
rect 22198 35334 22212 35386
rect 22236 35334 22250 35386
rect 22250 35334 22262 35386
rect 22262 35334 22292 35386
rect 22316 35334 22326 35386
rect 22326 35334 22372 35386
rect 22076 35332 22132 35334
rect 22156 35332 22212 35334
rect 22236 35332 22292 35334
rect 22316 35332 22372 35334
rect 22076 34298 22132 34300
rect 22156 34298 22212 34300
rect 22236 34298 22292 34300
rect 22316 34298 22372 34300
rect 22076 34246 22122 34298
rect 22122 34246 22132 34298
rect 22156 34246 22186 34298
rect 22186 34246 22198 34298
rect 22198 34246 22212 34298
rect 22236 34246 22250 34298
rect 22250 34246 22262 34298
rect 22262 34246 22292 34298
rect 22316 34246 22326 34298
rect 22326 34246 22372 34298
rect 22076 34244 22132 34246
rect 22156 34244 22212 34246
rect 22236 34244 22292 34246
rect 22316 34244 22372 34246
rect 22076 33210 22132 33212
rect 22156 33210 22212 33212
rect 22236 33210 22292 33212
rect 22316 33210 22372 33212
rect 22076 33158 22122 33210
rect 22122 33158 22132 33210
rect 22156 33158 22186 33210
rect 22186 33158 22198 33210
rect 22198 33158 22212 33210
rect 22236 33158 22250 33210
rect 22250 33158 22262 33210
rect 22262 33158 22292 33210
rect 22316 33158 22326 33210
rect 22326 33158 22372 33210
rect 22076 33156 22132 33158
rect 22156 33156 22212 33158
rect 22236 33156 22292 33158
rect 22316 33156 22372 33158
rect 22076 32122 22132 32124
rect 22156 32122 22212 32124
rect 22236 32122 22292 32124
rect 22316 32122 22372 32124
rect 22076 32070 22122 32122
rect 22122 32070 22132 32122
rect 22156 32070 22186 32122
rect 22186 32070 22198 32122
rect 22198 32070 22212 32122
rect 22236 32070 22250 32122
rect 22250 32070 22262 32122
rect 22262 32070 22292 32122
rect 22316 32070 22326 32122
rect 22326 32070 22372 32122
rect 22076 32068 22132 32070
rect 22156 32068 22212 32070
rect 22236 32068 22292 32070
rect 22316 32068 22372 32070
rect 13628 19066 13684 19068
rect 13708 19066 13764 19068
rect 13788 19066 13844 19068
rect 13868 19066 13924 19068
rect 13628 19014 13674 19066
rect 13674 19014 13684 19066
rect 13708 19014 13738 19066
rect 13738 19014 13750 19066
rect 13750 19014 13764 19066
rect 13788 19014 13802 19066
rect 13802 19014 13814 19066
rect 13814 19014 13844 19066
rect 13868 19014 13878 19066
rect 13878 19014 13924 19066
rect 13628 19012 13684 19014
rect 13708 19012 13764 19014
rect 13788 19012 13844 19014
rect 13868 19012 13924 19014
rect 13628 17978 13684 17980
rect 13708 17978 13764 17980
rect 13788 17978 13844 17980
rect 13868 17978 13924 17980
rect 13628 17926 13674 17978
rect 13674 17926 13684 17978
rect 13708 17926 13738 17978
rect 13738 17926 13750 17978
rect 13750 17926 13764 17978
rect 13788 17926 13802 17978
rect 13802 17926 13814 17978
rect 13814 17926 13844 17978
rect 13868 17926 13878 17978
rect 13878 17926 13924 17978
rect 13628 17924 13684 17926
rect 13708 17924 13764 17926
rect 13788 17924 13844 17926
rect 13868 17924 13924 17926
rect 13628 16890 13684 16892
rect 13708 16890 13764 16892
rect 13788 16890 13844 16892
rect 13868 16890 13924 16892
rect 13628 16838 13674 16890
rect 13674 16838 13684 16890
rect 13708 16838 13738 16890
rect 13738 16838 13750 16890
rect 13750 16838 13764 16890
rect 13788 16838 13802 16890
rect 13802 16838 13814 16890
rect 13814 16838 13844 16890
rect 13868 16838 13878 16890
rect 13878 16838 13924 16890
rect 13628 16836 13684 16838
rect 13708 16836 13764 16838
rect 13788 16836 13844 16838
rect 13868 16836 13924 16838
rect 13628 15802 13684 15804
rect 13708 15802 13764 15804
rect 13788 15802 13844 15804
rect 13868 15802 13924 15804
rect 13628 15750 13674 15802
rect 13674 15750 13684 15802
rect 13708 15750 13738 15802
rect 13738 15750 13750 15802
rect 13750 15750 13764 15802
rect 13788 15750 13802 15802
rect 13802 15750 13814 15802
rect 13814 15750 13844 15802
rect 13868 15750 13878 15802
rect 13878 15750 13924 15802
rect 13628 15748 13684 15750
rect 13708 15748 13764 15750
rect 13788 15748 13844 15750
rect 13868 15748 13924 15750
rect 13628 14714 13684 14716
rect 13708 14714 13764 14716
rect 13788 14714 13844 14716
rect 13868 14714 13924 14716
rect 13628 14662 13674 14714
rect 13674 14662 13684 14714
rect 13708 14662 13738 14714
rect 13738 14662 13750 14714
rect 13750 14662 13764 14714
rect 13788 14662 13802 14714
rect 13802 14662 13814 14714
rect 13814 14662 13844 14714
rect 13868 14662 13878 14714
rect 13878 14662 13924 14714
rect 13628 14660 13684 14662
rect 13708 14660 13764 14662
rect 13788 14660 13844 14662
rect 13868 14660 13924 14662
rect 13628 13626 13684 13628
rect 13708 13626 13764 13628
rect 13788 13626 13844 13628
rect 13868 13626 13924 13628
rect 13628 13574 13674 13626
rect 13674 13574 13684 13626
rect 13708 13574 13738 13626
rect 13738 13574 13750 13626
rect 13750 13574 13764 13626
rect 13788 13574 13802 13626
rect 13802 13574 13814 13626
rect 13814 13574 13844 13626
rect 13868 13574 13878 13626
rect 13878 13574 13924 13626
rect 13628 13572 13684 13574
rect 13708 13572 13764 13574
rect 13788 13572 13844 13574
rect 13868 13572 13924 13574
rect 13628 12538 13684 12540
rect 13708 12538 13764 12540
rect 13788 12538 13844 12540
rect 13868 12538 13924 12540
rect 13628 12486 13674 12538
rect 13674 12486 13684 12538
rect 13708 12486 13738 12538
rect 13738 12486 13750 12538
rect 13750 12486 13764 12538
rect 13788 12486 13802 12538
rect 13802 12486 13814 12538
rect 13814 12486 13844 12538
rect 13868 12486 13878 12538
rect 13878 12486 13924 12538
rect 13628 12484 13684 12486
rect 13708 12484 13764 12486
rect 13788 12484 13844 12486
rect 13868 12484 13924 12486
rect 13628 11450 13684 11452
rect 13708 11450 13764 11452
rect 13788 11450 13844 11452
rect 13868 11450 13924 11452
rect 13628 11398 13674 11450
rect 13674 11398 13684 11450
rect 13708 11398 13738 11450
rect 13738 11398 13750 11450
rect 13750 11398 13764 11450
rect 13788 11398 13802 11450
rect 13802 11398 13814 11450
rect 13814 11398 13844 11450
rect 13868 11398 13878 11450
rect 13878 11398 13924 11450
rect 13628 11396 13684 11398
rect 13708 11396 13764 11398
rect 13788 11396 13844 11398
rect 13868 11396 13924 11398
rect 13628 10362 13684 10364
rect 13708 10362 13764 10364
rect 13788 10362 13844 10364
rect 13868 10362 13924 10364
rect 13628 10310 13674 10362
rect 13674 10310 13684 10362
rect 13708 10310 13738 10362
rect 13738 10310 13750 10362
rect 13750 10310 13764 10362
rect 13788 10310 13802 10362
rect 13802 10310 13814 10362
rect 13814 10310 13844 10362
rect 13868 10310 13878 10362
rect 13878 10310 13924 10362
rect 13628 10308 13684 10310
rect 13708 10308 13764 10310
rect 13788 10308 13844 10310
rect 13868 10308 13924 10310
rect 13628 9274 13684 9276
rect 13708 9274 13764 9276
rect 13788 9274 13844 9276
rect 13868 9274 13924 9276
rect 13628 9222 13674 9274
rect 13674 9222 13684 9274
rect 13708 9222 13738 9274
rect 13738 9222 13750 9274
rect 13750 9222 13764 9274
rect 13788 9222 13802 9274
rect 13802 9222 13814 9274
rect 13814 9222 13844 9274
rect 13868 9222 13878 9274
rect 13878 9222 13924 9274
rect 13628 9220 13684 9222
rect 13708 9220 13764 9222
rect 13788 9220 13844 9222
rect 13868 9220 13924 9222
rect 13628 8186 13684 8188
rect 13708 8186 13764 8188
rect 13788 8186 13844 8188
rect 13868 8186 13924 8188
rect 13628 8134 13674 8186
rect 13674 8134 13684 8186
rect 13708 8134 13738 8186
rect 13738 8134 13750 8186
rect 13750 8134 13764 8186
rect 13788 8134 13802 8186
rect 13802 8134 13814 8186
rect 13814 8134 13844 8186
rect 13868 8134 13878 8186
rect 13878 8134 13924 8186
rect 13628 8132 13684 8134
rect 13708 8132 13764 8134
rect 13788 8132 13844 8134
rect 13868 8132 13924 8134
rect 13628 7098 13684 7100
rect 13708 7098 13764 7100
rect 13788 7098 13844 7100
rect 13868 7098 13924 7100
rect 13628 7046 13674 7098
rect 13674 7046 13684 7098
rect 13708 7046 13738 7098
rect 13738 7046 13750 7098
rect 13750 7046 13764 7098
rect 13788 7046 13802 7098
rect 13802 7046 13814 7098
rect 13814 7046 13844 7098
rect 13868 7046 13878 7098
rect 13878 7046 13924 7098
rect 13628 7044 13684 7046
rect 13708 7044 13764 7046
rect 13788 7044 13844 7046
rect 13868 7044 13924 7046
rect 13628 6010 13684 6012
rect 13708 6010 13764 6012
rect 13788 6010 13844 6012
rect 13868 6010 13924 6012
rect 13628 5958 13674 6010
rect 13674 5958 13684 6010
rect 13708 5958 13738 6010
rect 13738 5958 13750 6010
rect 13750 5958 13764 6010
rect 13788 5958 13802 6010
rect 13802 5958 13814 6010
rect 13814 5958 13844 6010
rect 13868 5958 13878 6010
rect 13878 5958 13924 6010
rect 13628 5956 13684 5958
rect 13708 5956 13764 5958
rect 13788 5956 13844 5958
rect 13868 5956 13924 5958
rect 13628 4922 13684 4924
rect 13708 4922 13764 4924
rect 13788 4922 13844 4924
rect 13868 4922 13924 4924
rect 13628 4870 13674 4922
rect 13674 4870 13684 4922
rect 13708 4870 13738 4922
rect 13738 4870 13750 4922
rect 13750 4870 13764 4922
rect 13788 4870 13802 4922
rect 13802 4870 13814 4922
rect 13814 4870 13844 4922
rect 13868 4870 13878 4922
rect 13878 4870 13924 4922
rect 13628 4868 13684 4870
rect 13708 4868 13764 4870
rect 13788 4868 13844 4870
rect 13868 4868 13924 4870
rect 13628 3834 13684 3836
rect 13708 3834 13764 3836
rect 13788 3834 13844 3836
rect 13868 3834 13924 3836
rect 13628 3782 13674 3834
rect 13674 3782 13684 3834
rect 13708 3782 13738 3834
rect 13738 3782 13750 3834
rect 13750 3782 13764 3834
rect 13788 3782 13802 3834
rect 13802 3782 13814 3834
rect 13814 3782 13844 3834
rect 13868 3782 13878 3834
rect 13878 3782 13924 3834
rect 13628 3780 13684 3782
rect 13708 3780 13764 3782
rect 13788 3780 13844 3782
rect 13868 3780 13924 3782
rect 13628 2746 13684 2748
rect 13708 2746 13764 2748
rect 13788 2746 13844 2748
rect 13868 2746 13924 2748
rect 13628 2694 13674 2746
rect 13674 2694 13684 2746
rect 13708 2694 13738 2746
rect 13738 2694 13750 2746
rect 13750 2694 13764 2746
rect 13788 2694 13802 2746
rect 13802 2694 13814 2746
rect 13814 2694 13844 2746
rect 13868 2694 13878 2746
rect 13878 2694 13924 2746
rect 13628 2692 13684 2694
rect 13708 2692 13764 2694
rect 13788 2692 13844 2694
rect 13868 2692 13924 2694
rect 17852 31578 17908 31580
rect 17932 31578 17988 31580
rect 18012 31578 18068 31580
rect 18092 31578 18148 31580
rect 17852 31526 17898 31578
rect 17898 31526 17908 31578
rect 17932 31526 17962 31578
rect 17962 31526 17974 31578
rect 17974 31526 17988 31578
rect 18012 31526 18026 31578
rect 18026 31526 18038 31578
rect 18038 31526 18068 31578
rect 18092 31526 18102 31578
rect 18102 31526 18148 31578
rect 17852 31524 17908 31526
rect 17932 31524 17988 31526
rect 18012 31524 18068 31526
rect 18092 31524 18148 31526
rect 17852 30490 17908 30492
rect 17932 30490 17988 30492
rect 18012 30490 18068 30492
rect 18092 30490 18148 30492
rect 17852 30438 17898 30490
rect 17898 30438 17908 30490
rect 17932 30438 17962 30490
rect 17962 30438 17974 30490
rect 17974 30438 17988 30490
rect 18012 30438 18026 30490
rect 18026 30438 18038 30490
rect 18038 30438 18068 30490
rect 18092 30438 18102 30490
rect 18102 30438 18148 30490
rect 17852 30436 17908 30438
rect 17932 30436 17988 30438
rect 18012 30436 18068 30438
rect 18092 30436 18148 30438
rect 17852 29402 17908 29404
rect 17932 29402 17988 29404
rect 18012 29402 18068 29404
rect 18092 29402 18148 29404
rect 17852 29350 17898 29402
rect 17898 29350 17908 29402
rect 17932 29350 17962 29402
rect 17962 29350 17974 29402
rect 17974 29350 17988 29402
rect 18012 29350 18026 29402
rect 18026 29350 18038 29402
rect 18038 29350 18068 29402
rect 18092 29350 18102 29402
rect 18102 29350 18148 29402
rect 17852 29348 17908 29350
rect 17932 29348 17988 29350
rect 18012 29348 18068 29350
rect 18092 29348 18148 29350
rect 17852 28314 17908 28316
rect 17932 28314 17988 28316
rect 18012 28314 18068 28316
rect 18092 28314 18148 28316
rect 17852 28262 17898 28314
rect 17898 28262 17908 28314
rect 17932 28262 17962 28314
rect 17962 28262 17974 28314
rect 17974 28262 17988 28314
rect 18012 28262 18026 28314
rect 18026 28262 18038 28314
rect 18038 28262 18068 28314
rect 18092 28262 18102 28314
rect 18102 28262 18148 28314
rect 17852 28260 17908 28262
rect 17932 28260 17988 28262
rect 18012 28260 18068 28262
rect 18092 28260 18148 28262
rect 17852 27226 17908 27228
rect 17932 27226 17988 27228
rect 18012 27226 18068 27228
rect 18092 27226 18148 27228
rect 17852 27174 17898 27226
rect 17898 27174 17908 27226
rect 17932 27174 17962 27226
rect 17962 27174 17974 27226
rect 17974 27174 17988 27226
rect 18012 27174 18026 27226
rect 18026 27174 18038 27226
rect 18038 27174 18068 27226
rect 18092 27174 18102 27226
rect 18102 27174 18148 27226
rect 17852 27172 17908 27174
rect 17932 27172 17988 27174
rect 18012 27172 18068 27174
rect 18092 27172 18148 27174
rect 17852 26138 17908 26140
rect 17932 26138 17988 26140
rect 18012 26138 18068 26140
rect 18092 26138 18148 26140
rect 17852 26086 17898 26138
rect 17898 26086 17908 26138
rect 17932 26086 17962 26138
rect 17962 26086 17974 26138
rect 17974 26086 17988 26138
rect 18012 26086 18026 26138
rect 18026 26086 18038 26138
rect 18038 26086 18068 26138
rect 18092 26086 18102 26138
rect 18102 26086 18148 26138
rect 17852 26084 17908 26086
rect 17932 26084 17988 26086
rect 18012 26084 18068 26086
rect 18092 26084 18148 26086
rect 17852 25050 17908 25052
rect 17932 25050 17988 25052
rect 18012 25050 18068 25052
rect 18092 25050 18148 25052
rect 17852 24998 17898 25050
rect 17898 24998 17908 25050
rect 17932 24998 17962 25050
rect 17962 24998 17974 25050
rect 17974 24998 17988 25050
rect 18012 24998 18026 25050
rect 18026 24998 18038 25050
rect 18038 24998 18068 25050
rect 18092 24998 18102 25050
rect 18102 24998 18148 25050
rect 17852 24996 17908 24998
rect 17932 24996 17988 24998
rect 18012 24996 18068 24998
rect 18092 24996 18148 24998
rect 17852 23962 17908 23964
rect 17932 23962 17988 23964
rect 18012 23962 18068 23964
rect 18092 23962 18148 23964
rect 17852 23910 17898 23962
rect 17898 23910 17908 23962
rect 17932 23910 17962 23962
rect 17962 23910 17974 23962
rect 17974 23910 17988 23962
rect 18012 23910 18026 23962
rect 18026 23910 18038 23962
rect 18038 23910 18068 23962
rect 18092 23910 18102 23962
rect 18102 23910 18148 23962
rect 17852 23908 17908 23910
rect 17932 23908 17988 23910
rect 18012 23908 18068 23910
rect 18092 23908 18148 23910
rect 17852 22874 17908 22876
rect 17932 22874 17988 22876
rect 18012 22874 18068 22876
rect 18092 22874 18148 22876
rect 17852 22822 17898 22874
rect 17898 22822 17908 22874
rect 17932 22822 17962 22874
rect 17962 22822 17974 22874
rect 17974 22822 17988 22874
rect 18012 22822 18026 22874
rect 18026 22822 18038 22874
rect 18038 22822 18068 22874
rect 18092 22822 18102 22874
rect 18102 22822 18148 22874
rect 17852 22820 17908 22822
rect 17932 22820 17988 22822
rect 18012 22820 18068 22822
rect 18092 22820 18148 22822
rect 17852 21786 17908 21788
rect 17932 21786 17988 21788
rect 18012 21786 18068 21788
rect 18092 21786 18148 21788
rect 17852 21734 17898 21786
rect 17898 21734 17908 21786
rect 17932 21734 17962 21786
rect 17962 21734 17974 21786
rect 17974 21734 17988 21786
rect 18012 21734 18026 21786
rect 18026 21734 18038 21786
rect 18038 21734 18068 21786
rect 18092 21734 18102 21786
rect 18102 21734 18148 21786
rect 17852 21732 17908 21734
rect 17932 21732 17988 21734
rect 18012 21732 18068 21734
rect 18092 21732 18148 21734
rect 17852 20698 17908 20700
rect 17932 20698 17988 20700
rect 18012 20698 18068 20700
rect 18092 20698 18148 20700
rect 17852 20646 17898 20698
rect 17898 20646 17908 20698
rect 17932 20646 17962 20698
rect 17962 20646 17974 20698
rect 17974 20646 17988 20698
rect 18012 20646 18026 20698
rect 18026 20646 18038 20698
rect 18038 20646 18068 20698
rect 18092 20646 18102 20698
rect 18102 20646 18148 20698
rect 17852 20644 17908 20646
rect 17932 20644 17988 20646
rect 18012 20644 18068 20646
rect 18092 20644 18148 20646
rect 17852 19610 17908 19612
rect 17932 19610 17988 19612
rect 18012 19610 18068 19612
rect 18092 19610 18148 19612
rect 17852 19558 17898 19610
rect 17898 19558 17908 19610
rect 17932 19558 17962 19610
rect 17962 19558 17974 19610
rect 17974 19558 17988 19610
rect 18012 19558 18026 19610
rect 18026 19558 18038 19610
rect 18038 19558 18068 19610
rect 18092 19558 18102 19610
rect 18102 19558 18148 19610
rect 17852 19556 17908 19558
rect 17932 19556 17988 19558
rect 18012 19556 18068 19558
rect 18092 19556 18148 19558
rect 22076 31034 22132 31036
rect 22156 31034 22212 31036
rect 22236 31034 22292 31036
rect 22316 31034 22372 31036
rect 22076 30982 22122 31034
rect 22122 30982 22132 31034
rect 22156 30982 22186 31034
rect 22186 30982 22198 31034
rect 22198 30982 22212 31034
rect 22236 30982 22250 31034
rect 22250 30982 22262 31034
rect 22262 30982 22292 31034
rect 22316 30982 22326 31034
rect 22326 30982 22372 31034
rect 22076 30980 22132 30982
rect 22156 30980 22212 30982
rect 22236 30980 22292 30982
rect 22316 30980 22372 30982
rect 17852 18522 17908 18524
rect 17932 18522 17988 18524
rect 18012 18522 18068 18524
rect 18092 18522 18148 18524
rect 17852 18470 17898 18522
rect 17898 18470 17908 18522
rect 17932 18470 17962 18522
rect 17962 18470 17974 18522
rect 17974 18470 17988 18522
rect 18012 18470 18026 18522
rect 18026 18470 18038 18522
rect 18038 18470 18068 18522
rect 18092 18470 18102 18522
rect 18102 18470 18148 18522
rect 17852 18468 17908 18470
rect 17932 18468 17988 18470
rect 18012 18468 18068 18470
rect 18092 18468 18148 18470
rect 17852 17434 17908 17436
rect 17932 17434 17988 17436
rect 18012 17434 18068 17436
rect 18092 17434 18148 17436
rect 17852 17382 17898 17434
rect 17898 17382 17908 17434
rect 17932 17382 17962 17434
rect 17962 17382 17974 17434
rect 17974 17382 17988 17434
rect 18012 17382 18026 17434
rect 18026 17382 18038 17434
rect 18038 17382 18068 17434
rect 18092 17382 18102 17434
rect 18102 17382 18148 17434
rect 17852 17380 17908 17382
rect 17932 17380 17988 17382
rect 18012 17380 18068 17382
rect 18092 17380 18148 17382
rect 17852 16346 17908 16348
rect 17932 16346 17988 16348
rect 18012 16346 18068 16348
rect 18092 16346 18148 16348
rect 17852 16294 17898 16346
rect 17898 16294 17908 16346
rect 17932 16294 17962 16346
rect 17962 16294 17974 16346
rect 17974 16294 17988 16346
rect 18012 16294 18026 16346
rect 18026 16294 18038 16346
rect 18038 16294 18068 16346
rect 18092 16294 18102 16346
rect 18102 16294 18148 16346
rect 17852 16292 17908 16294
rect 17932 16292 17988 16294
rect 18012 16292 18068 16294
rect 18092 16292 18148 16294
rect 17852 15258 17908 15260
rect 17932 15258 17988 15260
rect 18012 15258 18068 15260
rect 18092 15258 18148 15260
rect 17852 15206 17898 15258
rect 17898 15206 17908 15258
rect 17932 15206 17962 15258
rect 17962 15206 17974 15258
rect 17974 15206 17988 15258
rect 18012 15206 18026 15258
rect 18026 15206 18038 15258
rect 18038 15206 18068 15258
rect 18092 15206 18102 15258
rect 18102 15206 18148 15258
rect 17852 15204 17908 15206
rect 17932 15204 17988 15206
rect 18012 15204 18068 15206
rect 18092 15204 18148 15206
rect 17852 14170 17908 14172
rect 17932 14170 17988 14172
rect 18012 14170 18068 14172
rect 18092 14170 18148 14172
rect 17852 14118 17898 14170
rect 17898 14118 17908 14170
rect 17932 14118 17962 14170
rect 17962 14118 17974 14170
rect 17974 14118 17988 14170
rect 18012 14118 18026 14170
rect 18026 14118 18038 14170
rect 18038 14118 18068 14170
rect 18092 14118 18102 14170
rect 18102 14118 18148 14170
rect 17852 14116 17908 14118
rect 17932 14116 17988 14118
rect 18012 14116 18068 14118
rect 18092 14116 18148 14118
rect 17852 13082 17908 13084
rect 17932 13082 17988 13084
rect 18012 13082 18068 13084
rect 18092 13082 18148 13084
rect 17852 13030 17898 13082
rect 17898 13030 17908 13082
rect 17932 13030 17962 13082
rect 17962 13030 17974 13082
rect 17974 13030 17988 13082
rect 18012 13030 18026 13082
rect 18026 13030 18038 13082
rect 18038 13030 18068 13082
rect 18092 13030 18102 13082
rect 18102 13030 18148 13082
rect 17852 13028 17908 13030
rect 17932 13028 17988 13030
rect 18012 13028 18068 13030
rect 18092 13028 18148 13030
rect 17852 11994 17908 11996
rect 17932 11994 17988 11996
rect 18012 11994 18068 11996
rect 18092 11994 18148 11996
rect 17852 11942 17898 11994
rect 17898 11942 17908 11994
rect 17932 11942 17962 11994
rect 17962 11942 17974 11994
rect 17974 11942 17988 11994
rect 18012 11942 18026 11994
rect 18026 11942 18038 11994
rect 18038 11942 18068 11994
rect 18092 11942 18102 11994
rect 18102 11942 18148 11994
rect 17852 11940 17908 11942
rect 17932 11940 17988 11942
rect 18012 11940 18068 11942
rect 18092 11940 18148 11942
rect 17852 10906 17908 10908
rect 17932 10906 17988 10908
rect 18012 10906 18068 10908
rect 18092 10906 18148 10908
rect 17852 10854 17898 10906
rect 17898 10854 17908 10906
rect 17932 10854 17962 10906
rect 17962 10854 17974 10906
rect 17974 10854 17988 10906
rect 18012 10854 18026 10906
rect 18026 10854 18038 10906
rect 18038 10854 18068 10906
rect 18092 10854 18102 10906
rect 18102 10854 18148 10906
rect 17852 10852 17908 10854
rect 17932 10852 17988 10854
rect 18012 10852 18068 10854
rect 18092 10852 18148 10854
rect 17852 9818 17908 9820
rect 17932 9818 17988 9820
rect 18012 9818 18068 9820
rect 18092 9818 18148 9820
rect 17852 9766 17898 9818
rect 17898 9766 17908 9818
rect 17932 9766 17962 9818
rect 17962 9766 17974 9818
rect 17974 9766 17988 9818
rect 18012 9766 18026 9818
rect 18026 9766 18038 9818
rect 18038 9766 18068 9818
rect 18092 9766 18102 9818
rect 18102 9766 18148 9818
rect 17852 9764 17908 9766
rect 17932 9764 17988 9766
rect 18012 9764 18068 9766
rect 18092 9764 18148 9766
rect 17852 8730 17908 8732
rect 17932 8730 17988 8732
rect 18012 8730 18068 8732
rect 18092 8730 18148 8732
rect 17852 8678 17898 8730
rect 17898 8678 17908 8730
rect 17932 8678 17962 8730
rect 17962 8678 17974 8730
rect 17974 8678 17988 8730
rect 18012 8678 18026 8730
rect 18026 8678 18038 8730
rect 18038 8678 18068 8730
rect 18092 8678 18102 8730
rect 18102 8678 18148 8730
rect 17852 8676 17908 8678
rect 17932 8676 17988 8678
rect 18012 8676 18068 8678
rect 18092 8676 18148 8678
rect 17852 7642 17908 7644
rect 17932 7642 17988 7644
rect 18012 7642 18068 7644
rect 18092 7642 18148 7644
rect 17852 7590 17898 7642
rect 17898 7590 17908 7642
rect 17932 7590 17962 7642
rect 17962 7590 17974 7642
rect 17974 7590 17988 7642
rect 18012 7590 18026 7642
rect 18026 7590 18038 7642
rect 18038 7590 18068 7642
rect 18092 7590 18102 7642
rect 18102 7590 18148 7642
rect 17852 7588 17908 7590
rect 17932 7588 17988 7590
rect 18012 7588 18068 7590
rect 18092 7588 18148 7590
rect 17852 6554 17908 6556
rect 17932 6554 17988 6556
rect 18012 6554 18068 6556
rect 18092 6554 18148 6556
rect 17852 6502 17898 6554
rect 17898 6502 17908 6554
rect 17932 6502 17962 6554
rect 17962 6502 17974 6554
rect 17974 6502 17988 6554
rect 18012 6502 18026 6554
rect 18026 6502 18038 6554
rect 18038 6502 18068 6554
rect 18092 6502 18102 6554
rect 18102 6502 18148 6554
rect 17852 6500 17908 6502
rect 17932 6500 17988 6502
rect 18012 6500 18068 6502
rect 18092 6500 18148 6502
rect 22076 29946 22132 29948
rect 22156 29946 22212 29948
rect 22236 29946 22292 29948
rect 22316 29946 22372 29948
rect 22076 29894 22122 29946
rect 22122 29894 22132 29946
rect 22156 29894 22186 29946
rect 22186 29894 22198 29946
rect 22198 29894 22212 29946
rect 22236 29894 22250 29946
rect 22250 29894 22262 29946
rect 22262 29894 22292 29946
rect 22316 29894 22326 29946
rect 22326 29894 22372 29946
rect 22076 29892 22132 29894
rect 22156 29892 22212 29894
rect 22236 29892 22292 29894
rect 22316 29892 22372 29894
rect 22076 28858 22132 28860
rect 22156 28858 22212 28860
rect 22236 28858 22292 28860
rect 22316 28858 22372 28860
rect 22076 28806 22122 28858
rect 22122 28806 22132 28858
rect 22156 28806 22186 28858
rect 22186 28806 22198 28858
rect 22198 28806 22212 28858
rect 22236 28806 22250 28858
rect 22250 28806 22262 28858
rect 22262 28806 22292 28858
rect 22316 28806 22326 28858
rect 22326 28806 22372 28858
rect 22076 28804 22132 28806
rect 22156 28804 22212 28806
rect 22236 28804 22292 28806
rect 22316 28804 22372 28806
rect 22076 27770 22132 27772
rect 22156 27770 22212 27772
rect 22236 27770 22292 27772
rect 22316 27770 22372 27772
rect 22076 27718 22122 27770
rect 22122 27718 22132 27770
rect 22156 27718 22186 27770
rect 22186 27718 22198 27770
rect 22198 27718 22212 27770
rect 22236 27718 22250 27770
rect 22250 27718 22262 27770
rect 22262 27718 22292 27770
rect 22316 27718 22326 27770
rect 22326 27718 22372 27770
rect 22076 27716 22132 27718
rect 22156 27716 22212 27718
rect 22236 27716 22292 27718
rect 22316 27716 22372 27718
rect 22076 26682 22132 26684
rect 22156 26682 22212 26684
rect 22236 26682 22292 26684
rect 22316 26682 22372 26684
rect 22076 26630 22122 26682
rect 22122 26630 22132 26682
rect 22156 26630 22186 26682
rect 22186 26630 22198 26682
rect 22198 26630 22212 26682
rect 22236 26630 22250 26682
rect 22250 26630 22262 26682
rect 22262 26630 22292 26682
rect 22316 26630 22326 26682
rect 22326 26630 22372 26682
rect 22076 26628 22132 26630
rect 22156 26628 22212 26630
rect 22236 26628 22292 26630
rect 22316 26628 22372 26630
rect 22076 25594 22132 25596
rect 22156 25594 22212 25596
rect 22236 25594 22292 25596
rect 22316 25594 22372 25596
rect 22076 25542 22122 25594
rect 22122 25542 22132 25594
rect 22156 25542 22186 25594
rect 22186 25542 22198 25594
rect 22198 25542 22212 25594
rect 22236 25542 22250 25594
rect 22250 25542 22262 25594
rect 22262 25542 22292 25594
rect 22316 25542 22326 25594
rect 22326 25542 22372 25594
rect 22076 25540 22132 25542
rect 22156 25540 22212 25542
rect 22236 25540 22292 25542
rect 22316 25540 22372 25542
rect 22076 24506 22132 24508
rect 22156 24506 22212 24508
rect 22236 24506 22292 24508
rect 22316 24506 22372 24508
rect 22076 24454 22122 24506
rect 22122 24454 22132 24506
rect 22156 24454 22186 24506
rect 22186 24454 22198 24506
rect 22198 24454 22212 24506
rect 22236 24454 22250 24506
rect 22250 24454 22262 24506
rect 22262 24454 22292 24506
rect 22316 24454 22326 24506
rect 22326 24454 22372 24506
rect 22076 24452 22132 24454
rect 22156 24452 22212 24454
rect 22236 24452 22292 24454
rect 22316 24452 22372 24454
rect 22076 23418 22132 23420
rect 22156 23418 22212 23420
rect 22236 23418 22292 23420
rect 22316 23418 22372 23420
rect 22076 23366 22122 23418
rect 22122 23366 22132 23418
rect 22156 23366 22186 23418
rect 22186 23366 22198 23418
rect 22198 23366 22212 23418
rect 22236 23366 22250 23418
rect 22250 23366 22262 23418
rect 22262 23366 22292 23418
rect 22316 23366 22326 23418
rect 22326 23366 22372 23418
rect 22076 23364 22132 23366
rect 22156 23364 22212 23366
rect 22236 23364 22292 23366
rect 22316 23364 22372 23366
rect 22076 22330 22132 22332
rect 22156 22330 22212 22332
rect 22236 22330 22292 22332
rect 22316 22330 22372 22332
rect 22076 22278 22122 22330
rect 22122 22278 22132 22330
rect 22156 22278 22186 22330
rect 22186 22278 22198 22330
rect 22198 22278 22212 22330
rect 22236 22278 22250 22330
rect 22250 22278 22262 22330
rect 22262 22278 22292 22330
rect 22316 22278 22326 22330
rect 22326 22278 22372 22330
rect 22076 22276 22132 22278
rect 22156 22276 22212 22278
rect 22236 22276 22292 22278
rect 22316 22276 22372 22278
rect 26300 39194 26356 39196
rect 26380 39194 26436 39196
rect 26460 39194 26516 39196
rect 26540 39194 26596 39196
rect 26300 39142 26346 39194
rect 26346 39142 26356 39194
rect 26380 39142 26410 39194
rect 26410 39142 26422 39194
rect 26422 39142 26436 39194
rect 26460 39142 26474 39194
rect 26474 39142 26486 39194
rect 26486 39142 26516 39194
rect 26540 39142 26550 39194
rect 26550 39142 26596 39194
rect 26300 39140 26356 39142
rect 26380 39140 26436 39142
rect 26460 39140 26516 39142
rect 26540 39140 26596 39142
rect 26300 38106 26356 38108
rect 26380 38106 26436 38108
rect 26460 38106 26516 38108
rect 26540 38106 26596 38108
rect 26300 38054 26346 38106
rect 26346 38054 26356 38106
rect 26380 38054 26410 38106
rect 26410 38054 26422 38106
rect 26422 38054 26436 38106
rect 26460 38054 26474 38106
rect 26474 38054 26486 38106
rect 26486 38054 26516 38106
rect 26540 38054 26550 38106
rect 26550 38054 26596 38106
rect 26300 38052 26356 38054
rect 26380 38052 26436 38054
rect 26460 38052 26516 38054
rect 26540 38052 26596 38054
rect 26300 37018 26356 37020
rect 26380 37018 26436 37020
rect 26460 37018 26516 37020
rect 26540 37018 26596 37020
rect 26300 36966 26346 37018
rect 26346 36966 26356 37018
rect 26380 36966 26410 37018
rect 26410 36966 26422 37018
rect 26422 36966 26436 37018
rect 26460 36966 26474 37018
rect 26474 36966 26486 37018
rect 26486 36966 26516 37018
rect 26540 36966 26550 37018
rect 26550 36966 26596 37018
rect 26300 36964 26356 36966
rect 26380 36964 26436 36966
rect 26460 36964 26516 36966
rect 26540 36964 26596 36966
rect 26300 35930 26356 35932
rect 26380 35930 26436 35932
rect 26460 35930 26516 35932
rect 26540 35930 26596 35932
rect 26300 35878 26346 35930
rect 26346 35878 26356 35930
rect 26380 35878 26410 35930
rect 26410 35878 26422 35930
rect 26422 35878 26436 35930
rect 26460 35878 26474 35930
rect 26474 35878 26486 35930
rect 26486 35878 26516 35930
rect 26540 35878 26550 35930
rect 26550 35878 26596 35930
rect 26300 35876 26356 35878
rect 26380 35876 26436 35878
rect 26460 35876 26516 35878
rect 26540 35876 26596 35878
rect 26300 34842 26356 34844
rect 26380 34842 26436 34844
rect 26460 34842 26516 34844
rect 26540 34842 26596 34844
rect 26300 34790 26346 34842
rect 26346 34790 26356 34842
rect 26380 34790 26410 34842
rect 26410 34790 26422 34842
rect 26422 34790 26436 34842
rect 26460 34790 26474 34842
rect 26474 34790 26486 34842
rect 26486 34790 26516 34842
rect 26540 34790 26550 34842
rect 26550 34790 26596 34842
rect 26300 34788 26356 34790
rect 26380 34788 26436 34790
rect 26460 34788 26516 34790
rect 26540 34788 26596 34790
rect 26300 33754 26356 33756
rect 26380 33754 26436 33756
rect 26460 33754 26516 33756
rect 26540 33754 26596 33756
rect 26300 33702 26346 33754
rect 26346 33702 26356 33754
rect 26380 33702 26410 33754
rect 26410 33702 26422 33754
rect 26422 33702 26436 33754
rect 26460 33702 26474 33754
rect 26474 33702 26486 33754
rect 26486 33702 26516 33754
rect 26540 33702 26550 33754
rect 26550 33702 26596 33754
rect 26300 33700 26356 33702
rect 26380 33700 26436 33702
rect 26460 33700 26516 33702
rect 26540 33700 26596 33702
rect 26300 32666 26356 32668
rect 26380 32666 26436 32668
rect 26460 32666 26516 32668
rect 26540 32666 26596 32668
rect 26300 32614 26346 32666
rect 26346 32614 26356 32666
rect 26380 32614 26410 32666
rect 26410 32614 26422 32666
rect 26422 32614 26436 32666
rect 26460 32614 26474 32666
rect 26474 32614 26486 32666
rect 26486 32614 26516 32666
rect 26540 32614 26550 32666
rect 26550 32614 26596 32666
rect 26300 32612 26356 32614
rect 26380 32612 26436 32614
rect 26460 32612 26516 32614
rect 26540 32612 26596 32614
rect 26300 31578 26356 31580
rect 26380 31578 26436 31580
rect 26460 31578 26516 31580
rect 26540 31578 26596 31580
rect 26300 31526 26346 31578
rect 26346 31526 26356 31578
rect 26380 31526 26410 31578
rect 26410 31526 26422 31578
rect 26422 31526 26436 31578
rect 26460 31526 26474 31578
rect 26474 31526 26486 31578
rect 26486 31526 26516 31578
rect 26540 31526 26550 31578
rect 26550 31526 26596 31578
rect 26300 31524 26356 31526
rect 26380 31524 26436 31526
rect 26460 31524 26516 31526
rect 26540 31524 26596 31526
rect 31758 40840 31814 40896
rect 26300 30490 26356 30492
rect 26380 30490 26436 30492
rect 26460 30490 26516 30492
rect 26540 30490 26596 30492
rect 26300 30438 26346 30490
rect 26346 30438 26356 30490
rect 26380 30438 26410 30490
rect 26410 30438 26422 30490
rect 26422 30438 26436 30490
rect 26460 30438 26474 30490
rect 26474 30438 26486 30490
rect 26486 30438 26516 30490
rect 26540 30438 26550 30490
rect 26550 30438 26596 30490
rect 26300 30436 26356 30438
rect 26380 30436 26436 30438
rect 26460 30436 26516 30438
rect 26540 30436 26596 30438
rect 26300 29402 26356 29404
rect 26380 29402 26436 29404
rect 26460 29402 26516 29404
rect 26540 29402 26596 29404
rect 26300 29350 26346 29402
rect 26346 29350 26356 29402
rect 26380 29350 26410 29402
rect 26410 29350 26422 29402
rect 26422 29350 26436 29402
rect 26460 29350 26474 29402
rect 26474 29350 26486 29402
rect 26486 29350 26516 29402
rect 26540 29350 26550 29402
rect 26550 29350 26596 29402
rect 26300 29348 26356 29350
rect 26380 29348 26436 29350
rect 26460 29348 26516 29350
rect 26540 29348 26596 29350
rect 30524 39738 30580 39740
rect 30604 39738 30660 39740
rect 30684 39738 30740 39740
rect 30764 39738 30820 39740
rect 30524 39686 30570 39738
rect 30570 39686 30580 39738
rect 30604 39686 30634 39738
rect 30634 39686 30646 39738
rect 30646 39686 30660 39738
rect 30684 39686 30698 39738
rect 30698 39686 30710 39738
rect 30710 39686 30740 39738
rect 30764 39686 30774 39738
rect 30774 39686 30820 39738
rect 30524 39684 30580 39686
rect 30604 39684 30660 39686
rect 30684 39684 30740 39686
rect 30764 39684 30820 39686
rect 31758 38820 31814 38856
rect 31758 38800 31760 38820
rect 31760 38800 31812 38820
rect 31812 38800 31814 38820
rect 30524 38650 30580 38652
rect 30604 38650 30660 38652
rect 30684 38650 30740 38652
rect 30764 38650 30820 38652
rect 30524 38598 30570 38650
rect 30570 38598 30580 38650
rect 30604 38598 30634 38650
rect 30634 38598 30646 38650
rect 30646 38598 30660 38650
rect 30684 38598 30698 38650
rect 30698 38598 30710 38650
rect 30710 38598 30740 38650
rect 30764 38598 30774 38650
rect 30774 38598 30820 38650
rect 30524 38596 30580 38598
rect 30604 38596 30660 38598
rect 30684 38596 30740 38598
rect 30764 38596 30820 38598
rect 30524 37562 30580 37564
rect 30604 37562 30660 37564
rect 30684 37562 30740 37564
rect 30764 37562 30820 37564
rect 30524 37510 30570 37562
rect 30570 37510 30580 37562
rect 30604 37510 30634 37562
rect 30634 37510 30646 37562
rect 30646 37510 30660 37562
rect 30684 37510 30698 37562
rect 30698 37510 30710 37562
rect 30710 37510 30740 37562
rect 30764 37510 30774 37562
rect 30774 37510 30820 37562
rect 30524 37508 30580 37510
rect 30604 37508 30660 37510
rect 30684 37508 30740 37510
rect 30764 37508 30820 37510
rect 26300 28314 26356 28316
rect 26380 28314 26436 28316
rect 26460 28314 26516 28316
rect 26540 28314 26596 28316
rect 26300 28262 26346 28314
rect 26346 28262 26356 28314
rect 26380 28262 26410 28314
rect 26410 28262 26422 28314
rect 26422 28262 26436 28314
rect 26460 28262 26474 28314
rect 26474 28262 26486 28314
rect 26486 28262 26516 28314
rect 26540 28262 26550 28314
rect 26550 28262 26596 28314
rect 26300 28260 26356 28262
rect 26380 28260 26436 28262
rect 26460 28260 26516 28262
rect 26540 28260 26596 28262
rect 26300 27226 26356 27228
rect 26380 27226 26436 27228
rect 26460 27226 26516 27228
rect 26540 27226 26596 27228
rect 26300 27174 26346 27226
rect 26346 27174 26356 27226
rect 26380 27174 26410 27226
rect 26410 27174 26422 27226
rect 26422 27174 26436 27226
rect 26460 27174 26474 27226
rect 26474 27174 26486 27226
rect 26486 27174 26516 27226
rect 26540 27174 26550 27226
rect 26550 27174 26596 27226
rect 26300 27172 26356 27174
rect 26380 27172 26436 27174
rect 26460 27172 26516 27174
rect 26540 27172 26596 27174
rect 26300 26138 26356 26140
rect 26380 26138 26436 26140
rect 26460 26138 26516 26140
rect 26540 26138 26596 26140
rect 26300 26086 26346 26138
rect 26346 26086 26356 26138
rect 26380 26086 26410 26138
rect 26410 26086 26422 26138
rect 26422 26086 26436 26138
rect 26460 26086 26474 26138
rect 26474 26086 26486 26138
rect 26486 26086 26516 26138
rect 26540 26086 26550 26138
rect 26550 26086 26596 26138
rect 26300 26084 26356 26086
rect 26380 26084 26436 26086
rect 26460 26084 26516 26086
rect 26540 26084 26596 26086
rect 26300 25050 26356 25052
rect 26380 25050 26436 25052
rect 26460 25050 26516 25052
rect 26540 25050 26596 25052
rect 26300 24998 26346 25050
rect 26346 24998 26356 25050
rect 26380 24998 26410 25050
rect 26410 24998 26422 25050
rect 26422 24998 26436 25050
rect 26460 24998 26474 25050
rect 26474 24998 26486 25050
rect 26486 24998 26516 25050
rect 26540 24998 26550 25050
rect 26550 24998 26596 25050
rect 26300 24996 26356 24998
rect 26380 24996 26436 24998
rect 26460 24996 26516 24998
rect 26540 24996 26596 24998
rect 26300 23962 26356 23964
rect 26380 23962 26436 23964
rect 26460 23962 26516 23964
rect 26540 23962 26596 23964
rect 26300 23910 26346 23962
rect 26346 23910 26356 23962
rect 26380 23910 26410 23962
rect 26410 23910 26422 23962
rect 26422 23910 26436 23962
rect 26460 23910 26474 23962
rect 26474 23910 26486 23962
rect 26486 23910 26516 23962
rect 26540 23910 26550 23962
rect 26550 23910 26596 23962
rect 26300 23908 26356 23910
rect 26380 23908 26436 23910
rect 26460 23908 26516 23910
rect 26540 23908 26596 23910
rect 26300 22874 26356 22876
rect 26380 22874 26436 22876
rect 26460 22874 26516 22876
rect 26540 22874 26596 22876
rect 26300 22822 26346 22874
rect 26346 22822 26356 22874
rect 26380 22822 26410 22874
rect 26410 22822 26422 22874
rect 26422 22822 26436 22874
rect 26460 22822 26474 22874
rect 26474 22822 26486 22874
rect 26486 22822 26516 22874
rect 26540 22822 26550 22874
rect 26550 22822 26596 22874
rect 26300 22820 26356 22822
rect 26380 22820 26436 22822
rect 26460 22820 26516 22822
rect 26540 22820 26596 22822
rect 26300 21786 26356 21788
rect 26380 21786 26436 21788
rect 26460 21786 26516 21788
rect 26540 21786 26596 21788
rect 26300 21734 26346 21786
rect 26346 21734 26356 21786
rect 26380 21734 26410 21786
rect 26410 21734 26422 21786
rect 26422 21734 26436 21786
rect 26460 21734 26474 21786
rect 26474 21734 26486 21786
rect 26486 21734 26516 21786
rect 26540 21734 26550 21786
rect 26550 21734 26596 21786
rect 26300 21732 26356 21734
rect 26380 21732 26436 21734
rect 26460 21732 26516 21734
rect 26540 21732 26596 21734
rect 22076 21242 22132 21244
rect 22156 21242 22212 21244
rect 22236 21242 22292 21244
rect 22316 21242 22372 21244
rect 22076 21190 22122 21242
rect 22122 21190 22132 21242
rect 22156 21190 22186 21242
rect 22186 21190 22198 21242
rect 22198 21190 22212 21242
rect 22236 21190 22250 21242
rect 22250 21190 22262 21242
rect 22262 21190 22292 21242
rect 22316 21190 22326 21242
rect 22326 21190 22372 21242
rect 22076 21188 22132 21190
rect 22156 21188 22212 21190
rect 22236 21188 22292 21190
rect 22316 21188 22372 21190
rect 22076 20154 22132 20156
rect 22156 20154 22212 20156
rect 22236 20154 22292 20156
rect 22316 20154 22372 20156
rect 22076 20102 22122 20154
rect 22122 20102 22132 20154
rect 22156 20102 22186 20154
rect 22186 20102 22198 20154
rect 22198 20102 22212 20154
rect 22236 20102 22250 20154
rect 22250 20102 22262 20154
rect 22262 20102 22292 20154
rect 22316 20102 22326 20154
rect 22326 20102 22372 20154
rect 22076 20100 22132 20102
rect 22156 20100 22212 20102
rect 22236 20100 22292 20102
rect 22316 20100 22372 20102
rect 26300 20698 26356 20700
rect 26380 20698 26436 20700
rect 26460 20698 26516 20700
rect 26540 20698 26596 20700
rect 26300 20646 26346 20698
rect 26346 20646 26356 20698
rect 26380 20646 26410 20698
rect 26410 20646 26422 20698
rect 26422 20646 26436 20698
rect 26460 20646 26474 20698
rect 26474 20646 26486 20698
rect 26486 20646 26516 20698
rect 26540 20646 26550 20698
rect 26550 20646 26596 20698
rect 26300 20644 26356 20646
rect 26380 20644 26436 20646
rect 26460 20644 26516 20646
rect 26540 20644 26596 20646
rect 26300 19610 26356 19612
rect 26380 19610 26436 19612
rect 26460 19610 26516 19612
rect 26540 19610 26596 19612
rect 26300 19558 26346 19610
rect 26346 19558 26356 19610
rect 26380 19558 26410 19610
rect 26410 19558 26422 19610
rect 26422 19558 26436 19610
rect 26460 19558 26474 19610
rect 26474 19558 26486 19610
rect 26486 19558 26516 19610
rect 26540 19558 26550 19610
rect 26550 19558 26596 19610
rect 26300 19556 26356 19558
rect 26380 19556 26436 19558
rect 26460 19556 26516 19558
rect 26540 19556 26596 19558
rect 22076 19066 22132 19068
rect 22156 19066 22212 19068
rect 22236 19066 22292 19068
rect 22316 19066 22372 19068
rect 22076 19014 22122 19066
rect 22122 19014 22132 19066
rect 22156 19014 22186 19066
rect 22186 19014 22198 19066
rect 22198 19014 22212 19066
rect 22236 19014 22250 19066
rect 22250 19014 22262 19066
rect 22262 19014 22292 19066
rect 22316 19014 22326 19066
rect 22326 19014 22372 19066
rect 22076 19012 22132 19014
rect 22156 19012 22212 19014
rect 22236 19012 22292 19014
rect 22316 19012 22372 19014
rect 26300 18522 26356 18524
rect 26380 18522 26436 18524
rect 26460 18522 26516 18524
rect 26540 18522 26596 18524
rect 26300 18470 26346 18522
rect 26346 18470 26356 18522
rect 26380 18470 26410 18522
rect 26410 18470 26422 18522
rect 26422 18470 26436 18522
rect 26460 18470 26474 18522
rect 26474 18470 26486 18522
rect 26486 18470 26516 18522
rect 26540 18470 26550 18522
rect 26550 18470 26596 18522
rect 26300 18468 26356 18470
rect 26380 18468 26436 18470
rect 26460 18468 26516 18470
rect 26540 18468 26596 18470
rect 22076 17978 22132 17980
rect 22156 17978 22212 17980
rect 22236 17978 22292 17980
rect 22316 17978 22372 17980
rect 22076 17926 22122 17978
rect 22122 17926 22132 17978
rect 22156 17926 22186 17978
rect 22186 17926 22198 17978
rect 22198 17926 22212 17978
rect 22236 17926 22250 17978
rect 22250 17926 22262 17978
rect 22262 17926 22292 17978
rect 22316 17926 22326 17978
rect 22326 17926 22372 17978
rect 22076 17924 22132 17926
rect 22156 17924 22212 17926
rect 22236 17924 22292 17926
rect 22316 17924 22372 17926
rect 22076 16890 22132 16892
rect 22156 16890 22212 16892
rect 22236 16890 22292 16892
rect 22316 16890 22372 16892
rect 22076 16838 22122 16890
rect 22122 16838 22132 16890
rect 22156 16838 22186 16890
rect 22186 16838 22198 16890
rect 22198 16838 22212 16890
rect 22236 16838 22250 16890
rect 22250 16838 22262 16890
rect 22262 16838 22292 16890
rect 22316 16838 22326 16890
rect 22326 16838 22372 16890
rect 22076 16836 22132 16838
rect 22156 16836 22212 16838
rect 22236 16836 22292 16838
rect 22316 16836 22372 16838
rect 22076 15802 22132 15804
rect 22156 15802 22212 15804
rect 22236 15802 22292 15804
rect 22316 15802 22372 15804
rect 22076 15750 22122 15802
rect 22122 15750 22132 15802
rect 22156 15750 22186 15802
rect 22186 15750 22198 15802
rect 22198 15750 22212 15802
rect 22236 15750 22250 15802
rect 22250 15750 22262 15802
rect 22262 15750 22292 15802
rect 22316 15750 22326 15802
rect 22326 15750 22372 15802
rect 22076 15748 22132 15750
rect 22156 15748 22212 15750
rect 22236 15748 22292 15750
rect 22316 15748 22372 15750
rect 17852 5466 17908 5468
rect 17932 5466 17988 5468
rect 18012 5466 18068 5468
rect 18092 5466 18148 5468
rect 17852 5414 17898 5466
rect 17898 5414 17908 5466
rect 17932 5414 17962 5466
rect 17962 5414 17974 5466
rect 17974 5414 17988 5466
rect 18012 5414 18026 5466
rect 18026 5414 18038 5466
rect 18038 5414 18068 5466
rect 18092 5414 18102 5466
rect 18102 5414 18148 5466
rect 17852 5412 17908 5414
rect 17932 5412 17988 5414
rect 18012 5412 18068 5414
rect 18092 5412 18148 5414
rect 17852 4378 17908 4380
rect 17932 4378 17988 4380
rect 18012 4378 18068 4380
rect 18092 4378 18148 4380
rect 17852 4326 17898 4378
rect 17898 4326 17908 4378
rect 17932 4326 17962 4378
rect 17962 4326 17974 4378
rect 17974 4326 17988 4378
rect 18012 4326 18026 4378
rect 18026 4326 18038 4378
rect 18038 4326 18068 4378
rect 18092 4326 18102 4378
rect 18102 4326 18148 4378
rect 17852 4324 17908 4326
rect 17932 4324 17988 4326
rect 18012 4324 18068 4326
rect 18092 4324 18148 4326
rect 17852 3290 17908 3292
rect 17932 3290 17988 3292
rect 18012 3290 18068 3292
rect 18092 3290 18148 3292
rect 17852 3238 17898 3290
rect 17898 3238 17908 3290
rect 17932 3238 17962 3290
rect 17962 3238 17974 3290
rect 17974 3238 17988 3290
rect 18012 3238 18026 3290
rect 18026 3238 18038 3290
rect 18038 3238 18068 3290
rect 18092 3238 18102 3290
rect 18102 3238 18148 3290
rect 17852 3236 17908 3238
rect 17932 3236 17988 3238
rect 18012 3236 18068 3238
rect 18092 3236 18148 3238
rect 17852 2202 17908 2204
rect 17932 2202 17988 2204
rect 18012 2202 18068 2204
rect 18092 2202 18148 2204
rect 17852 2150 17898 2202
rect 17898 2150 17908 2202
rect 17932 2150 17962 2202
rect 17962 2150 17974 2202
rect 17974 2150 17988 2202
rect 18012 2150 18026 2202
rect 18026 2150 18038 2202
rect 18038 2150 18068 2202
rect 18092 2150 18102 2202
rect 18102 2150 18148 2202
rect 17852 2148 17908 2150
rect 17932 2148 17988 2150
rect 18012 2148 18068 2150
rect 18092 2148 18148 2150
rect 22076 14714 22132 14716
rect 22156 14714 22212 14716
rect 22236 14714 22292 14716
rect 22316 14714 22372 14716
rect 22076 14662 22122 14714
rect 22122 14662 22132 14714
rect 22156 14662 22186 14714
rect 22186 14662 22198 14714
rect 22198 14662 22212 14714
rect 22236 14662 22250 14714
rect 22250 14662 22262 14714
rect 22262 14662 22292 14714
rect 22316 14662 22326 14714
rect 22326 14662 22372 14714
rect 22076 14660 22132 14662
rect 22156 14660 22212 14662
rect 22236 14660 22292 14662
rect 22316 14660 22372 14662
rect 22076 13626 22132 13628
rect 22156 13626 22212 13628
rect 22236 13626 22292 13628
rect 22316 13626 22372 13628
rect 22076 13574 22122 13626
rect 22122 13574 22132 13626
rect 22156 13574 22186 13626
rect 22186 13574 22198 13626
rect 22198 13574 22212 13626
rect 22236 13574 22250 13626
rect 22250 13574 22262 13626
rect 22262 13574 22292 13626
rect 22316 13574 22326 13626
rect 22326 13574 22372 13626
rect 22076 13572 22132 13574
rect 22156 13572 22212 13574
rect 22236 13572 22292 13574
rect 22316 13572 22372 13574
rect 26300 17434 26356 17436
rect 26380 17434 26436 17436
rect 26460 17434 26516 17436
rect 26540 17434 26596 17436
rect 26300 17382 26346 17434
rect 26346 17382 26356 17434
rect 26380 17382 26410 17434
rect 26410 17382 26422 17434
rect 26422 17382 26436 17434
rect 26460 17382 26474 17434
rect 26474 17382 26486 17434
rect 26486 17382 26516 17434
rect 26540 17382 26550 17434
rect 26550 17382 26596 17434
rect 26300 17380 26356 17382
rect 26380 17380 26436 17382
rect 26460 17380 26516 17382
rect 26540 17380 26596 17382
rect 26300 16346 26356 16348
rect 26380 16346 26436 16348
rect 26460 16346 26516 16348
rect 26540 16346 26596 16348
rect 26300 16294 26346 16346
rect 26346 16294 26356 16346
rect 26380 16294 26410 16346
rect 26410 16294 26422 16346
rect 26422 16294 26436 16346
rect 26460 16294 26474 16346
rect 26474 16294 26486 16346
rect 26486 16294 26516 16346
rect 26540 16294 26550 16346
rect 26550 16294 26596 16346
rect 26300 16292 26356 16294
rect 26380 16292 26436 16294
rect 26460 16292 26516 16294
rect 26540 16292 26596 16294
rect 26300 15258 26356 15260
rect 26380 15258 26436 15260
rect 26460 15258 26516 15260
rect 26540 15258 26596 15260
rect 26300 15206 26346 15258
rect 26346 15206 26356 15258
rect 26380 15206 26410 15258
rect 26410 15206 26422 15258
rect 26422 15206 26436 15258
rect 26460 15206 26474 15258
rect 26474 15206 26486 15258
rect 26486 15206 26516 15258
rect 26540 15206 26550 15258
rect 26550 15206 26596 15258
rect 26300 15204 26356 15206
rect 26380 15204 26436 15206
rect 26460 15204 26516 15206
rect 26540 15204 26596 15206
rect 26300 14170 26356 14172
rect 26380 14170 26436 14172
rect 26460 14170 26516 14172
rect 26540 14170 26596 14172
rect 26300 14118 26346 14170
rect 26346 14118 26356 14170
rect 26380 14118 26410 14170
rect 26410 14118 26422 14170
rect 26422 14118 26436 14170
rect 26460 14118 26474 14170
rect 26474 14118 26486 14170
rect 26486 14118 26516 14170
rect 26540 14118 26550 14170
rect 26550 14118 26596 14170
rect 26300 14116 26356 14118
rect 26380 14116 26436 14118
rect 26460 14116 26516 14118
rect 26540 14116 26596 14118
rect 26300 13082 26356 13084
rect 26380 13082 26436 13084
rect 26460 13082 26516 13084
rect 26540 13082 26596 13084
rect 26300 13030 26346 13082
rect 26346 13030 26356 13082
rect 26380 13030 26410 13082
rect 26410 13030 26422 13082
rect 26422 13030 26436 13082
rect 26460 13030 26474 13082
rect 26474 13030 26486 13082
rect 26486 13030 26516 13082
rect 26540 13030 26550 13082
rect 26550 13030 26596 13082
rect 26300 13028 26356 13030
rect 26380 13028 26436 13030
rect 26460 13028 26516 13030
rect 26540 13028 26596 13030
rect 22076 12538 22132 12540
rect 22156 12538 22212 12540
rect 22236 12538 22292 12540
rect 22316 12538 22372 12540
rect 22076 12486 22122 12538
rect 22122 12486 22132 12538
rect 22156 12486 22186 12538
rect 22186 12486 22198 12538
rect 22198 12486 22212 12538
rect 22236 12486 22250 12538
rect 22250 12486 22262 12538
rect 22262 12486 22292 12538
rect 22316 12486 22326 12538
rect 22326 12486 22372 12538
rect 22076 12484 22132 12486
rect 22156 12484 22212 12486
rect 22236 12484 22292 12486
rect 22316 12484 22372 12486
rect 22076 11450 22132 11452
rect 22156 11450 22212 11452
rect 22236 11450 22292 11452
rect 22316 11450 22372 11452
rect 22076 11398 22122 11450
rect 22122 11398 22132 11450
rect 22156 11398 22186 11450
rect 22186 11398 22198 11450
rect 22198 11398 22212 11450
rect 22236 11398 22250 11450
rect 22250 11398 22262 11450
rect 22262 11398 22292 11450
rect 22316 11398 22326 11450
rect 22326 11398 22372 11450
rect 22076 11396 22132 11398
rect 22156 11396 22212 11398
rect 22236 11396 22292 11398
rect 22316 11396 22372 11398
rect 22076 10362 22132 10364
rect 22156 10362 22212 10364
rect 22236 10362 22292 10364
rect 22316 10362 22372 10364
rect 22076 10310 22122 10362
rect 22122 10310 22132 10362
rect 22156 10310 22186 10362
rect 22186 10310 22198 10362
rect 22198 10310 22212 10362
rect 22236 10310 22250 10362
rect 22250 10310 22262 10362
rect 22262 10310 22292 10362
rect 22316 10310 22326 10362
rect 22326 10310 22372 10362
rect 22076 10308 22132 10310
rect 22156 10308 22212 10310
rect 22236 10308 22292 10310
rect 22316 10308 22372 10310
rect 22076 9274 22132 9276
rect 22156 9274 22212 9276
rect 22236 9274 22292 9276
rect 22316 9274 22372 9276
rect 22076 9222 22122 9274
rect 22122 9222 22132 9274
rect 22156 9222 22186 9274
rect 22186 9222 22198 9274
rect 22198 9222 22212 9274
rect 22236 9222 22250 9274
rect 22250 9222 22262 9274
rect 22262 9222 22292 9274
rect 22316 9222 22326 9274
rect 22326 9222 22372 9274
rect 22076 9220 22132 9222
rect 22156 9220 22212 9222
rect 22236 9220 22292 9222
rect 22316 9220 22372 9222
rect 22076 8186 22132 8188
rect 22156 8186 22212 8188
rect 22236 8186 22292 8188
rect 22316 8186 22372 8188
rect 22076 8134 22122 8186
rect 22122 8134 22132 8186
rect 22156 8134 22186 8186
rect 22186 8134 22198 8186
rect 22198 8134 22212 8186
rect 22236 8134 22250 8186
rect 22250 8134 22262 8186
rect 22262 8134 22292 8186
rect 22316 8134 22326 8186
rect 22326 8134 22372 8186
rect 22076 8132 22132 8134
rect 22156 8132 22212 8134
rect 22236 8132 22292 8134
rect 22316 8132 22372 8134
rect 22076 7098 22132 7100
rect 22156 7098 22212 7100
rect 22236 7098 22292 7100
rect 22316 7098 22372 7100
rect 22076 7046 22122 7098
rect 22122 7046 22132 7098
rect 22156 7046 22186 7098
rect 22186 7046 22198 7098
rect 22198 7046 22212 7098
rect 22236 7046 22250 7098
rect 22250 7046 22262 7098
rect 22262 7046 22292 7098
rect 22316 7046 22326 7098
rect 22326 7046 22372 7098
rect 22076 7044 22132 7046
rect 22156 7044 22212 7046
rect 22236 7044 22292 7046
rect 22316 7044 22372 7046
rect 22076 6010 22132 6012
rect 22156 6010 22212 6012
rect 22236 6010 22292 6012
rect 22316 6010 22372 6012
rect 22076 5958 22122 6010
rect 22122 5958 22132 6010
rect 22156 5958 22186 6010
rect 22186 5958 22198 6010
rect 22198 5958 22212 6010
rect 22236 5958 22250 6010
rect 22250 5958 22262 6010
rect 22262 5958 22292 6010
rect 22316 5958 22326 6010
rect 22326 5958 22372 6010
rect 22076 5956 22132 5958
rect 22156 5956 22212 5958
rect 22236 5956 22292 5958
rect 22316 5956 22372 5958
rect 22076 4922 22132 4924
rect 22156 4922 22212 4924
rect 22236 4922 22292 4924
rect 22316 4922 22372 4924
rect 22076 4870 22122 4922
rect 22122 4870 22132 4922
rect 22156 4870 22186 4922
rect 22186 4870 22198 4922
rect 22198 4870 22212 4922
rect 22236 4870 22250 4922
rect 22250 4870 22262 4922
rect 22262 4870 22292 4922
rect 22316 4870 22326 4922
rect 22326 4870 22372 4922
rect 22076 4868 22132 4870
rect 22156 4868 22212 4870
rect 22236 4868 22292 4870
rect 22316 4868 22372 4870
rect 22076 3834 22132 3836
rect 22156 3834 22212 3836
rect 22236 3834 22292 3836
rect 22316 3834 22372 3836
rect 22076 3782 22122 3834
rect 22122 3782 22132 3834
rect 22156 3782 22186 3834
rect 22186 3782 22198 3834
rect 22198 3782 22212 3834
rect 22236 3782 22250 3834
rect 22250 3782 22262 3834
rect 22262 3782 22292 3834
rect 22316 3782 22326 3834
rect 22326 3782 22372 3834
rect 22076 3780 22132 3782
rect 22156 3780 22212 3782
rect 22236 3780 22292 3782
rect 22316 3780 22372 3782
rect 22076 2746 22132 2748
rect 22156 2746 22212 2748
rect 22236 2746 22292 2748
rect 22316 2746 22372 2748
rect 22076 2694 22122 2746
rect 22122 2694 22132 2746
rect 22156 2694 22186 2746
rect 22186 2694 22198 2746
rect 22198 2694 22212 2746
rect 22236 2694 22250 2746
rect 22250 2694 22262 2746
rect 22262 2694 22292 2746
rect 22316 2694 22326 2746
rect 22326 2694 22372 2746
rect 22076 2692 22132 2694
rect 22156 2692 22212 2694
rect 22236 2692 22292 2694
rect 22316 2692 22372 2694
rect 26300 11994 26356 11996
rect 26380 11994 26436 11996
rect 26460 11994 26516 11996
rect 26540 11994 26596 11996
rect 26300 11942 26346 11994
rect 26346 11942 26356 11994
rect 26380 11942 26410 11994
rect 26410 11942 26422 11994
rect 26422 11942 26436 11994
rect 26460 11942 26474 11994
rect 26474 11942 26486 11994
rect 26486 11942 26516 11994
rect 26540 11942 26550 11994
rect 26550 11942 26596 11994
rect 26300 11940 26356 11942
rect 26380 11940 26436 11942
rect 26460 11940 26516 11942
rect 26540 11940 26596 11942
rect 26300 10906 26356 10908
rect 26380 10906 26436 10908
rect 26460 10906 26516 10908
rect 26540 10906 26596 10908
rect 26300 10854 26346 10906
rect 26346 10854 26356 10906
rect 26380 10854 26410 10906
rect 26410 10854 26422 10906
rect 26422 10854 26436 10906
rect 26460 10854 26474 10906
rect 26474 10854 26486 10906
rect 26486 10854 26516 10906
rect 26540 10854 26550 10906
rect 26550 10854 26596 10906
rect 26300 10852 26356 10854
rect 26380 10852 26436 10854
rect 26460 10852 26516 10854
rect 26540 10852 26596 10854
rect 31666 36760 31722 36816
rect 30524 36474 30580 36476
rect 30604 36474 30660 36476
rect 30684 36474 30740 36476
rect 30764 36474 30820 36476
rect 30524 36422 30570 36474
rect 30570 36422 30580 36474
rect 30604 36422 30634 36474
rect 30634 36422 30646 36474
rect 30646 36422 30660 36474
rect 30684 36422 30698 36474
rect 30698 36422 30710 36474
rect 30710 36422 30740 36474
rect 30764 36422 30774 36474
rect 30774 36422 30820 36474
rect 30524 36420 30580 36422
rect 30604 36420 30660 36422
rect 30684 36420 30740 36422
rect 30764 36420 30820 36422
rect 30524 35386 30580 35388
rect 30604 35386 30660 35388
rect 30684 35386 30740 35388
rect 30764 35386 30820 35388
rect 30524 35334 30570 35386
rect 30570 35334 30580 35386
rect 30604 35334 30634 35386
rect 30634 35334 30646 35386
rect 30646 35334 30660 35386
rect 30684 35334 30698 35386
rect 30698 35334 30710 35386
rect 30710 35334 30740 35386
rect 30764 35334 30774 35386
rect 30774 35334 30820 35386
rect 30524 35332 30580 35334
rect 30604 35332 30660 35334
rect 30684 35332 30740 35334
rect 30764 35332 30820 35334
rect 31574 34720 31630 34776
rect 30524 34298 30580 34300
rect 30604 34298 30660 34300
rect 30684 34298 30740 34300
rect 30764 34298 30820 34300
rect 30524 34246 30570 34298
rect 30570 34246 30580 34298
rect 30604 34246 30634 34298
rect 30634 34246 30646 34298
rect 30646 34246 30660 34298
rect 30684 34246 30698 34298
rect 30698 34246 30710 34298
rect 30710 34246 30740 34298
rect 30764 34246 30774 34298
rect 30774 34246 30820 34298
rect 30524 34244 30580 34246
rect 30604 34244 30660 34246
rect 30684 34244 30740 34246
rect 30764 34244 30820 34246
rect 30524 33210 30580 33212
rect 30604 33210 30660 33212
rect 30684 33210 30740 33212
rect 30764 33210 30820 33212
rect 30524 33158 30570 33210
rect 30570 33158 30580 33210
rect 30604 33158 30634 33210
rect 30634 33158 30646 33210
rect 30646 33158 30660 33210
rect 30684 33158 30698 33210
rect 30698 33158 30710 33210
rect 30710 33158 30740 33210
rect 30764 33158 30774 33210
rect 30774 33158 30820 33210
rect 30524 33156 30580 33158
rect 30604 33156 30660 33158
rect 30684 33156 30740 33158
rect 30764 33156 30820 33158
rect 30524 32122 30580 32124
rect 30604 32122 30660 32124
rect 30684 32122 30740 32124
rect 30764 32122 30820 32124
rect 30524 32070 30570 32122
rect 30570 32070 30580 32122
rect 30604 32070 30634 32122
rect 30634 32070 30646 32122
rect 30646 32070 30660 32122
rect 30684 32070 30698 32122
rect 30698 32070 30710 32122
rect 30710 32070 30740 32122
rect 30764 32070 30774 32122
rect 30774 32070 30820 32122
rect 30524 32068 30580 32070
rect 30604 32068 30660 32070
rect 30684 32068 30740 32070
rect 30764 32068 30820 32070
rect 30524 31034 30580 31036
rect 30604 31034 30660 31036
rect 30684 31034 30740 31036
rect 30764 31034 30820 31036
rect 30524 30982 30570 31034
rect 30570 30982 30580 31034
rect 30604 30982 30634 31034
rect 30634 30982 30646 31034
rect 30646 30982 30660 31034
rect 30684 30982 30698 31034
rect 30698 30982 30710 31034
rect 30710 30982 30740 31034
rect 30764 30982 30774 31034
rect 30774 30982 30820 31034
rect 30524 30980 30580 30982
rect 30604 30980 30660 30982
rect 30684 30980 30740 30982
rect 30764 30980 30820 30982
rect 30524 29946 30580 29948
rect 30604 29946 30660 29948
rect 30684 29946 30740 29948
rect 30764 29946 30820 29948
rect 30524 29894 30570 29946
rect 30570 29894 30580 29946
rect 30604 29894 30634 29946
rect 30634 29894 30646 29946
rect 30646 29894 30660 29946
rect 30684 29894 30698 29946
rect 30698 29894 30710 29946
rect 30710 29894 30740 29946
rect 30764 29894 30774 29946
rect 30774 29894 30820 29946
rect 30524 29892 30580 29894
rect 30604 29892 30660 29894
rect 30684 29892 30740 29894
rect 30764 29892 30820 29894
rect 30524 28858 30580 28860
rect 30604 28858 30660 28860
rect 30684 28858 30740 28860
rect 30764 28858 30820 28860
rect 30524 28806 30570 28858
rect 30570 28806 30580 28858
rect 30604 28806 30634 28858
rect 30634 28806 30646 28858
rect 30646 28806 30660 28858
rect 30684 28806 30698 28858
rect 30698 28806 30710 28858
rect 30710 28806 30740 28858
rect 30764 28806 30774 28858
rect 30774 28806 30820 28858
rect 30524 28804 30580 28806
rect 30604 28804 30660 28806
rect 30684 28804 30740 28806
rect 30764 28804 30820 28806
rect 32586 39480 32642 39536
rect 32310 33396 32312 33416
rect 32312 33396 32364 33416
rect 32364 33396 32366 33416
rect 32310 33360 32366 33396
rect 30524 27770 30580 27772
rect 30604 27770 30660 27772
rect 30684 27770 30740 27772
rect 30764 27770 30820 27772
rect 30524 27718 30570 27770
rect 30570 27718 30580 27770
rect 30604 27718 30634 27770
rect 30634 27718 30646 27770
rect 30646 27718 30660 27770
rect 30684 27718 30698 27770
rect 30698 27718 30710 27770
rect 30710 27718 30740 27770
rect 30764 27718 30774 27770
rect 30774 27718 30820 27770
rect 30524 27716 30580 27718
rect 30604 27716 30660 27718
rect 30684 27716 30740 27718
rect 30764 27716 30820 27718
rect 30524 26682 30580 26684
rect 30604 26682 30660 26684
rect 30684 26682 30740 26684
rect 30764 26682 30820 26684
rect 30524 26630 30570 26682
rect 30570 26630 30580 26682
rect 30604 26630 30634 26682
rect 30634 26630 30646 26682
rect 30646 26630 30660 26682
rect 30684 26630 30698 26682
rect 30698 26630 30710 26682
rect 30710 26630 30740 26682
rect 30764 26630 30774 26682
rect 30774 26630 30820 26682
rect 30524 26628 30580 26630
rect 30604 26628 30660 26630
rect 30684 26628 30740 26630
rect 30764 26628 30820 26630
rect 30524 25594 30580 25596
rect 30604 25594 30660 25596
rect 30684 25594 30740 25596
rect 30764 25594 30820 25596
rect 30524 25542 30570 25594
rect 30570 25542 30580 25594
rect 30604 25542 30634 25594
rect 30634 25542 30646 25594
rect 30646 25542 30660 25594
rect 30684 25542 30698 25594
rect 30698 25542 30710 25594
rect 30710 25542 30740 25594
rect 30764 25542 30774 25594
rect 30774 25542 30820 25594
rect 30524 25540 30580 25542
rect 30604 25540 30660 25542
rect 30684 25540 30740 25542
rect 30764 25540 30820 25542
rect 31758 25200 31814 25256
rect 30524 24506 30580 24508
rect 30604 24506 30660 24508
rect 30684 24506 30740 24508
rect 30764 24506 30820 24508
rect 30524 24454 30570 24506
rect 30570 24454 30580 24506
rect 30604 24454 30634 24506
rect 30634 24454 30646 24506
rect 30646 24454 30660 24506
rect 30684 24454 30698 24506
rect 30698 24454 30710 24506
rect 30710 24454 30740 24506
rect 30764 24454 30774 24506
rect 30774 24454 30820 24506
rect 30524 24452 30580 24454
rect 30604 24452 30660 24454
rect 30684 24452 30740 24454
rect 30764 24452 30820 24454
rect 30524 23418 30580 23420
rect 30604 23418 30660 23420
rect 30684 23418 30740 23420
rect 30764 23418 30820 23420
rect 30524 23366 30570 23418
rect 30570 23366 30580 23418
rect 30604 23366 30634 23418
rect 30634 23366 30646 23418
rect 30646 23366 30660 23418
rect 30684 23366 30698 23418
rect 30698 23366 30710 23418
rect 30710 23366 30740 23418
rect 30764 23366 30774 23418
rect 30774 23366 30820 23418
rect 30524 23364 30580 23366
rect 30604 23364 30660 23366
rect 30684 23364 30740 23366
rect 30764 23364 30820 23366
rect 30524 22330 30580 22332
rect 30604 22330 30660 22332
rect 30684 22330 30740 22332
rect 30764 22330 30820 22332
rect 30524 22278 30570 22330
rect 30570 22278 30580 22330
rect 30604 22278 30634 22330
rect 30634 22278 30646 22330
rect 30646 22278 30660 22330
rect 30684 22278 30698 22330
rect 30698 22278 30710 22330
rect 30710 22278 30740 22330
rect 30764 22278 30774 22330
rect 30774 22278 30820 22330
rect 30524 22276 30580 22278
rect 30604 22276 30660 22278
rect 30684 22276 30740 22278
rect 30764 22276 30820 22278
rect 30524 21242 30580 21244
rect 30604 21242 30660 21244
rect 30684 21242 30740 21244
rect 30764 21242 30820 21244
rect 30524 21190 30570 21242
rect 30570 21190 30580 21242
rect 30604 21190 30634 21242
rect 30634 21190 30646 21242
rect 30646 21190 30660 21242
rect 30684 21190 30698 21242
rect 30698 21190 30710 21242
rect 30710 21190 30740 21242
rect 30764 21190 30774 21242
rect 30774 21190 30820 21242
rect 30524 21188 30580 21190
rect 30604 21188 30660 21190
rect 30684 21188 30740 21190
rect 30764 21188 30820 21190
rect 30524 20154 30580 20156
rect 30604 20154 30660 20156
rect 30684 20154 30740 20156
rect 30764 20154 30820 20156
rect 30524 20102 30570 20154
rect 30570 20102 30580 20154
rect 30604 20102 30634 20154
rect 30634 20102 30646 20154
rect 30646 20102 30660 20154
rect 30684 20102 30698 20154
rect 30698 20102 30710 20154
rect 30710 20102 30740 20154
rect 30764 20102 30774 20154
rect 30774 20102 30820 20154
rect 30524 20100 30580 20102
rect 30604 20100 30660 20102
rect 30684 20100 30740 20102
rect 30764 20100 30820 20102
rect 26300 9818 26356 9820
rect 26380 9818 26436 9820
rect 26460 9818 26516 9820
rect 26540 9818 26596 9820
rect 26300 9766 26346 9818
rect 26346 9766 26356 9818
rect 26380 9766 26410 9818
rect 26410 9766 26422 9818
rect 26422 9766 26436 9818
rect 26460 9766 26474 9818
rect 26474 9766 26486 9818
rect 26486 9766 26516 9818
rect 26540 9766 26550 9818
rect 26550 9766 26596 9818
rect 26300 9764 26356 9766
rect 26380 9764 26436 9766
rect 26460 9764 26516 9766
rect 26540 9764 26596 9766
rect 26300 8730 26356 8732
rect 26380 8730 26436 8732
rect 26460 8730 26516 8732
rect 26540 8730 26596 8732
rect 26300 8678 26346 8730
rect 26346 8678 26356 8730
rect 26380 8678 26410 8730
rect 26410 8678 26422 8730
rect 26422 8678 26436 8730
rect 26460 8678 26474 8730
rect 26474 8678 26486 8730
rect 26486 8678 26516 8730
rect 26540 8678 26550 8730
rect 26550 8678 26596 8730
rect 26300 8676 26356 8678
rect 26380 8676 26436 8678
rect 26460 8676 26516 8678
rect 26540 8676 26596 8678
rect 26300 7642 26356 7644
rect 26380 7642 26436 7644
rect 26460 7642 26516 7644
rect 26540 7642 26596 7644
rect 26300 7590 26346 7642
rect 26346 7590 26356 7642
rect 26380 7590 26410 7642
rect 26410 7590 26422 7642
rect 26422 7590 26436 7642
rect 26460 7590 26474 7642
rect 26474 7590 26486 7642
rect 26486 7590 26516 7642
rect 26540 7590 26550 7642
rect 26550 7590 26596 7642
rect 26300 7588 26356 7590
rect 26380 7588 26436 7590
rect 26460 7588 26516 7590
rect 26540 7588 26596 7590
rect 26300 6554 26356 6556
rect 26380 6554 26436 6556
rect 26460 6554 26516 6556
rect 26540 6554 26596 6556
rect 26300 6502 26346 6554
rect 26346 6502 26356 6554
rect 26380 6502 26410 6554
rect 26410 6502 26422 6554
rect 26422 6502 26436 6554
rect 26460 6502 26474 6554
rect 26474 6502 26486 6554
rect 26486 6502 26516 6554
rect 26540 6502 26550 6554
rect 26550 6502 26596 6554
rect 26300 6500 26356 6502
rect 26380 6500 26436 6502
rect 26460 6500 26516 6502
rect 26540 6500 26596 6502
rect 26300 5466 26356 5468
rect 26380 5466 26436 5468
rect 26460 5466 26516 5468
rect 26540 5466 26596 5468
rect 26300 5414 26346 5466
rect 26346 5414 26356 5466
rect 26380 5414 26410 5466
rect 26410 5414 26422 5466
rect 26422 5414 26436 5466
rect 26460 5414 26474 5466
rect 26474 5414 26486 5466
rect 26486 5414 26516 5466
rect 26540 5414 26550 5466
rect 26550 5414 26596 5466
rect 26300 5412 26356 5414
rect 26380 5412 26436 5414
rect 26460 5412 26516 5414
rect 26540 5412 26596 5414
rect 26300 4378 26356 4380
rect 26380 4378 26436 4380
rect 26460 4378 26516 4380
rect 26540 4378 26596 4380
rect 26300 4326 26346 4378
rect 26346 4326 26356 4378
rect 26380 4326 26410 4378
rect 26410 4326 26422 4378
rect 26422 4326 26436 4378
rect 26460 4326 26474 4378
rect 26474 4326 26486 4378
rect 26486 4326 26516 4378
rect 26540 4326 26550 4378
rect 26550 4326 26596 4378
rect 26300 4324 26356 4326
rect 26380 4324 26436 4326
rect 26460 4324 26516 4326
rect 26540 4324 26596 4326
rect 26300 3290 26356 3292
rect 26380 3290 26436 3292
rect 26460 3290 26516 3292
rect 26540 3290 26596 3292
rect 26300 3238 26346 3290
rect 26346 3238 26356 3290
rect 26380 3238 26410 3290
rect 26410 3238 26422 3290
rect 26422 3238 26436 3290
rect 26460 3238 26474 3290
rect 26474 3238 26486 3290
rect 26486 3238 26516 3290
rect 26540 3238 26550 3290
rect 26550 3238 26596 3290
rect 26300 3236 26356 3238
rect 26380 3236 26436 3238
rect 26460 3236 26516 3238
rect 26540 3236 26596 3238
rect 26300 2202 26356 2204
rect 26380 2202 26436 2204
rect 26460 2202 26516 2204
rect 26540 2202 26596 2204
rect 26300 2150 26346 2202
rect 26346 2150 26356 2202
rect 26380 2150 26410 2202
rect 26410 2150 26422 2202
rect 26422 2150 26436 2202
rect 26460 2150 26474 2202
rect 26474 2150 26486 2202
rect 26486 2150 26516 2202
rect 26540 2150 26550 2202
rect 26550 2150 26596 2202
rect 26300 2148 26356 2150
rect 26380 2148 26436 2150
rect 26460 2148 26516 2150
rect 26540 2148 26596 2150
rect 30524 19066 30580 19068
rect 30604 19066 30660 19068
rect 30684 19066 30740 19068
rect 30764 19066 30820 19068
rect 30524 19014 30570 19066
rect 30570 19014 30580 19066
rect 30604 19014 30634 19066
rect 30634 19014 30646 19066
rect 30646 19014 30660 19066
rect 30684 19014 30698 19066
rect 30698 19014 30710 19066
rect 30710 19014 30740 19066
rect 30764 19014 30774 19066
rect 30774 19014 30820 19066
rect 30524 19012 30580 19014
rect 30604 19012 30660 19014
rect 30684 19012 30740 19014
rect 30764 19012 30820 19014
rect 30524 17978 30580 17980
rect 30604 17978 30660 17980
rect 30684 17978 30740 17980
rect 30764 17978 30820 17980
rect 30524 17926 30570 17978
rect 30570 17926 30580 17978
rect 30604 17926 30634 17978
rect 30634 17926 30646 17978
rect 30646 17926 30660 17978
rect 30684 17926 30698 17978
rect 30698 17926 30710 17978
rect 30710 17926 30740 17978
rect 30764 17926 30774 17978
rect 30774 17926 30820 17978
rect 30524 17924 30580 17926
rect 30604 17924 30660 17926
rect 30684 17924 30740 17926
rect 30764 17924 30820 17926
rect 30524 16890 30580 16892
rect 30604 16890 30660 16892
rect 30684 16890 30740 16892
rect 30764 16890 30820 16892
rect 30524 16838 30570 16890
rect 30570 16838 30580 16890
rect 30604 16838 30634 16890
rect 30634 16838 30646 16890
rect 30646 16838 30660 16890
rect 30684 16838 30698 16890
rect 30698 16838 30710 16890
rect 30710 16838 30740 16890
rect 30764 16838 30774 16890
rect 30774 16838 30820 16890
rect 30524 16836 30580 16838
rect 30604 16836 30660 16838
rect 30684 16836 30740 16838
rect 30764 16836 30820 16838
rect 30524 15802 30580 15804
rect 30604 15802 30660 15804
rect 30684 15802 30740 15804
rect 30764 15802 30820 15804
rect 30524 15750 30570 15802
rect 30570 15750 30580 15802
rect 30604 15750 30634 15802
rect 30634 15750 30646 15802
rect 30646 15750 30660 15802
rect 30684 15750 30698 15802
rect 30698 15750 30710 15802
rect 30710 15750 30740 15802
rect 30764 15750 30774 15802
rect 30774 15750 30820 15802
rect 30524 15748 30580 15750
rect 30604 15748 30660 15750
rect 30684 15748 30740 15750
rect 30764 15748 30820 15750
rect 30524 14714 30580 14716
rect 30604 14714 30660 14716
rect 30684 14714 30740 14716
rect 30764 14714 30820 14716
rect 30524 14662 30570 14714
rect 30570 14662 30580 14714
rect 30604 14662 30634 14714
rect 30634 14662 30646 14714
rect 30646 14662 30660 14714
rect 30684 14662 30698 14714
rect 30698 14662 30710 14714
rect 30710 14662 30740 14714
rect 30764 14662 30774 14714
rect 30774 14662 30820 14714
rect 30524 14660 30580 14662
rect 30604 14660 30660 14662
rect 30684 14660 30740 14662
rect 30764 14660 30820 14662
rect 30524 13626 30580 13628
rect 30604 13626 30660 13628
rect 30684 13626 30740 13628
rect 30764 13626 30820 13628
rect 30524 13574 30570 13626
rect 30570 13574 30580 13626
rect 30604 13574 30634 13626
rect 30634 13574 30646 13626
rect 30646 13574 30660 13626
rect 30684 13574 30698 13626
rect 30698 13574 30710 13626
rect 30710 13574 30740 13626
rect 30764 13574 30774 13626
rect 30774 13574 30820 13626
rect 30524 13572 30580 13574
rect 30604 13572 30660 13574
rect 30684 13572 30740 13574
rect 30764 13572 30820 13574
rect 30524 12538 30580 12540
rect 30604 12538 30660 12540
rect 30684 12538 30740 12540
rect 30764 12538 30820 12540
rect 30524 12486 30570 12538
rect 30570 12486 30580 12538
rect 30604 12486 30634 12538
rect 30634 12486 30646 12538
rect 30646 12486 30660 12538
rect 30684 12486 30698 12538
rect 30698 12486 30710 12538
rect 30710 12486 30740 12538
rect 30764 12486 30774 12538
rect 30774 12486 30820 12538
rect 30524 12484 30580 12486
rect 30604 12484 30660 12486
rect 30684 12484 30740 12486
rect 30764 12484 30820 12486
rect 30524 11450 30580 11452
rect 30604 11450 30660 11452
rect 30684 11450 30740 11452
rect 30764 11450 30820 11452
rect 30524 11398 30570 11450
rect 30570 11398 30580 11450
rect 30604 11398 30634 11450
rect 30634 11398 30646 11450
rect 30646 11398 30660 11450
rect 30684 11398 30698 11450
rect 30698 11398 30710 11450
rect 30710 11398 30740 11450
rect 30764 11398 30774 11450
rect 30774 11398 30820 11450
rect 30524 11396 30580 11398
rect 30604 11396 30660 11398
rect 30684 11396 30740 11398
rect 30764 11396 30820 11398
rect 30524 10362 30580 10364
rect 30604 10362 30660 10364
rect 30684 10362 30740 10364
rect 30764 10362 30820 10364
rect 30524 10310 30570 10362
rect 30570 10310 30580 10362
rect 30604 10310 30634 10362
rect 30634 10310 30646 10362
rect 30646 10310 30660 10362
rect 30684 10310 30698 10362
rect 30698 10310 30710 10362
rect 30710 10310 30740 10362
rect 30764 10310 30774 10362
rect 30774 10310 30820 10362
rect 30524 10308 30580 10310
rect 30604 10308 30660 10310
rect 30684 10308 30740 10310
rect 30764 10308 30820 10310
rect 30524 9274 30580 9276
rect 30604 9274 30660 9276
rect 30684 9274 30740 9276
rect 30764 9274 30820 9276
rect 30524 9222 30570 9274
rect 30570 9222 30580 9274
rect 30604 9222 30634 9274
rect 30634 9222 30646 9274
rect 30646 9222 30660 9274
rect 30684 9222 30698 9274
rect 30698 9222 30710 9274
rect 30710 9222 30740 9274
rect 30764 9222 30774 9274
rect 30774 9222 30820 9274
rect 30524 9220 30580 9222
rect 30604 9220 30660 9222
rect 30684 9220 30740 9222
rect 30764 9220 30820 9222
rect 30524 8186 30580 8188
rect 30604 8186 30660 8188
rect 30684 8186 30740 8188
rect 30764 8186 30820 8188
rect 30524 8134 30570 8186
rect 30570 8134 30580 8186
rect 30604 8134 30634 8186
rect 30634 8134 30646 8186
rect 30646 8134 30660 8186
rect 30684 8134 30698 8186
rect 30698 8134 30710 8186
rect 30710 8134 30740 8186
rect 30764 8134 30774 8186
rect 30774 8134 30820 8186
rect 30524 8132 30580 8134
rect 30604 8132 30660 8134
rect 30684 8132 30740 8134
rect 30764 8132 30820 8134
rect 30524 7098 30580 7100
rect 30604 7098 30660 7100
rect 30684 7098 30740 7100
rect 30764 7098 30820 7100
rect 30524 7046 30570 7098
rect 30570 7046 30580 7098
rect 30604 7046 30634 7098
rect 30634 7046 30646 7098
rect 30646 7046 30660 7098
rect 30684 7046 30698 7098
rect 30698 7046 30710 7098
rect 30710 7046 30740 7098
rect 30764 7046 30774 7098
rect 30774 7046 30820 7098
rect 30524 7044 30580 7046
rect 30604 7044 30660 7046
rect 30684 7044 30740 7046
rect 30764 7044 30820 7046
rect 30524 6010 30580 6012
rect 30604 6010 30660 6012
rect 30684 6010 30740 6012
rect 30764 6010 30820 6012
rect 30524 5958 30570 6010
rect 30570 5958 30580 6010
rect 30604 5958 30634 6010
rect 30634 5958 30646 6010
rect 30646 5958 30660 6010
rect 30684 5958 30698 6010
rect 30698 5958 30710 6010
rect 30710 5958 30740 6010
rect 30764 5958 30774 6010
rect 30774 5958 30820 6010
rect 30524 5956 30580 5958
rect 30604 5956 30660 5958
rect 30684 5956 30740 5958
rect 30764 5956 30820 5958
rect 30524 4922 30580 4924
rect 30604 4922 30660 4924
rect 30684 4922 30740 4924
rect 30764 4922 30820 4924
rect 30524 4870 30570 4922
rect 30570 4870 30580 4922
rect 30604 4870 30634 4922
rect 30634 4870 30646 4922
rect 30646 4870 30660 4922
rect 30684 4870 30698 4922
rect 30698 4870 30710 4922
rect 30710 4870 30740 4922
rect 30764 4870 30774 4922
rect 30774 4870 30820 4922
rect 30524 4868 30580 4870
rect 30604 4868 30660 4870
rect 30684 4868 30740 4870
rect 30764 4868 30820 4870
rect 30524 3834 30580 3836
rect 30604 3834 30660 3836
rect 30684 3834 30740 3836
rect 30764 3834 30820 3836
rect 30524 3782 30570 3834
rect 30570 3782 30580 3834
rect 30604 3782 30634 3834
rect 30634 3782 30646 3834
rect 30646 3782 30660 3834
rect 30684 3782 30698 3834
rect 30698 3782 30710 3834
rect 30710 3782 30740 3834
rect 30764 3782 30774 3834
rect 30774 3782 30820 3834
rect 30524 3780 30580 3782
rect 30604 3780 30660 3782
rect 30684 3780 30740 3782
rect 30764 3780 30820 3782
rect 30524 2746 30580 2748
rect 30604 2746 30660 2748
rect 30684 2746 30740 2748
rect 30764 2746 30820 2748
rect 30524 2694 30570 2746
rect 30570 2694 30580 2746
rect 30604 2694 30634 2746
rect 30634 2694 30646 2746
rect 30646 2694 30660 2746
rect 30684 2694 30698 2746
rect 30698 2694 30710 2746
rect 30710 2694 30740 2746
rect 30764 2694 30774 2746
rect 30774 2694 30820 2746
rect 30524 2692 30580 2694
rect 30604 2692 30660 2694
rect 30684 2692 30740 2694
rect 30764 2692 30820 2694
rect 31758 19760 31814 19816
rect 32954 34040 33010 34096
rect 32310 17076 32312 17096
rect 32312 17076 32364 17096
rect 32364 17076 32366 17096
rect 32310 17040 32366 17076
rect 33046 32000 33102 32056
rect 34150 38120 34206 38176
rect 33690 32680 33746 32736
rect 34150 31320 34206 31376
rect 33046 27920 33102 27976
rect 33046 25916 33048 25936
rect 33048 25916 33100 25936
rect 33100 25916 33102 25936
rect 33046 25880 33102 25916
rect 32678 24520 32734 24576
rect 32954 20476 32956 20496
rect 32956 20476 33008 20496
rect 33008 20476 33010 20496
rect 32954 20440 33010 20476
rect 33046 19080 33102 19136
rect 33046 17740 33102 17776
rect 33046 17720 33048 17740
rect 33048 17720 33100 17740
rect 33100 17720 33102 17740
rect 34150 23840 34206 23896
rect 34150 23160 34206 23216
rect 31758 14340 31814 14376
rect 31758 14320 31760 14340
rect 31760 14320 31812 14340
rect 31812 14320 31814 14340
rect 32770 13640 32826 13696
rect 33046 12280 33102 12336
rect 31758 8880 31814 8936
rect 31758 2080 31814 2136
rect 32310 4800 32366 4856
rect 32402 4120 32458 4176
rect 34150 16360 34206 16416
rect 34150 12960 34206 13016
rect 33046 3440 33102 3496
rect 31390 720 31446 776
rect 34150 6860 34206 6896
rect 34150 6840 34152 6860
rect 34152 6840 34204 6860
rect 34204 6840 34206 6860
rect 33966 40 34022 96
<< metal3 >>
rect 0 41578 800 41668
rect 3601 41578 3667 41581
rect 0 41576 3667 41578
rect 0 41520 3606 41576
rect 3662 41520 3667 41576
rect 0 41518 3667 41520
rect 0 41428 800 41518
rect 3601 41515 3667 41518
rect 0 40898 800 40988
rect 4061 40898 4127 40901
rect 0 40896 4127 40898
rect 0 40840 4066 40896
rect 4122 40840 4127 40896
rect 0 40838 4127 40840
rect 0 40748 800 40838
rect 4061 40835 4127 40838
rect 31753 40898 31819 40901
rect 35200 40898 36000 40988
rect 31753 40896 36000 40898
rect 31753 40840 31758 40896
rect 31814 40840 36000 40896
rect 31753 40838 36000 40840
rect 31753 40835 31819 40838
rect 35200 40748 36000 40838
rect 35200 40068 36000 40308
rect 5170 39744 5486 39745
rect 5170 39680 5176 39744
rect 5240 39680 5256 39744
rect 5320 39680 5336 39744
rect 5400 39680 5416 39744
rect 5480 39680 5486 39744
rect 5170 39679 5486 39680
rect 13618 39744 13934 39745
rect 13618 39680 13624 39744
rect 13688 39680 13704 39744
rect 13768 39680 13784 39744
rect 13848 39680 13864 39744
rect 13928 39680 13934 39744
rect 13618 39679 13934 39680
rect 22066 39744 22382 39745
rect 22066 39680 22072 39744
rect 22136 39680 22152 39744
rect 22216 39680 22232 39744
rect 22296 39680 22312 39744
rect 22376 39680 22382 39744
rect 22066 39679 22382 39680
rect 30514 39744 30830 39745
rect 30514 39680 30520 39744
rect 30584 39680 30600 39744
rect 30664 39680 30680 39744
rect 30744 39680 30760 39744
rect 30824 39680 30830 39744
rect 30514 39679 30830 39680
rect 0 39388 800 39628
rect 32581 39538 32647 39541
rect 35200 39538 36000 39628
rect 32581 39536 36000 39538
rect 32581 39480 32586 39536
rect 32642 39480 36000 39536
rect 32581 39478 36000 39480
rect 32581 39475 32647 39478
rect 35200 39388 36000 39478
rect 9394 39200 9710 39201
rect 9394 39136 9400 39200
rect 9464 39136 9480 39200
rect 9544 39136 9560 39200
rect 9624 39136 9640 39200
rect 9704 39136 9710 39200
rect 9394 39135 9710 39136
rect 17842 39200 18158 39201
rect 17842 39136 17848 39200
rect 17912 39136 17928 39200
rect 17992 39136 18008 39200
rect 18072 39136 18088 39200
rect 18152 39136 18158 39200
rect 17842 39135 18158 39136
rect 26290 39200 26606 39201
rect 26290 39136 26296 39200
rect 26360 39136 26376 39200
rect 26440 39136 26456 39200
rect 26520 39136 26536 39200
rect 26600 39136 26606 39200
rect 26290 39135 26606 39136
rect 0 38708 800 38948
rect 31753 38858 31819 38861
rect 35200 38858 36000 38948
rect 31753 38856 36000 38858
rect 31753 38800 31758 38856
rect 31814 38800 36000 38856
rect 31753 38798 36000 38800
rect 31753 38795 31819 38798
rect 35200 38708 36000 38798
rect 5170 38656 5486 38657
rect 5170 38592 5176 38656
rect 5240 38592 5256 38656
rect 5320 38592 5336 38656
rect 5400 38592 5416 38656
rect 5480 38592 5486 38656
rect 5170 38591 5486 38592
rect 13618 38656 13934 38657
rect 13618 38592 13624 38656
rect 13688 38592 13704 38656
rect 13768 38592 13784 38656
rect 13848 38592 13864 38656
rect 13928 38592 13934 38656
rect 13618 38591 13934 38592
rect 22066 38656 22382 38657
rect 22066 38592 22072 38656
rect 22136 38592 22152 38656
rect 22216 38592 22232 38656
rect 22296 38592 22312 38656
rect 22376 38592 22382 38656
rect 22066 38591 22382 38592
rect 30514 38656 30830 38657
rect 30514 38592 30520 38656
rect 30584 38592 30600 38656
rect 30664 38592 30680 38656
rect 30744 38592 30760 38656
rect 30824 38592 30830 38656
rect 30514 38591 30830 38592
rect 0 38028 800 38268
rect 34145 38178 34211 38181
rect 35200 38178 36000 38268
rect 34145 38176 36000 38178
rect 34145 38120 34150 38176
rect 34206 38120 36000 38176
rect 34145 38118 36000 38120
rect 34145 38115 34211 38118
rect 9394 38112 9710 38113
rect 9394 38048 9400 38112
rect 9464 38048 9480 38112
rect 9544 38048 9560 38112
rect 9624 38048 9640 38112
rect 9704 38048 9710 38112
rect 9394 38047 9710 38048
rect 17842 38112 18158 38113
rect 17842 38048 17848 38112
rect 17912 38048 17928 38112
rect 17992 38048 18008 38112
rect 18072 38048 18088 38112
rect 18152 38048 18158 38112
rect 17842 38047 18158 38048
rect 26290 38112 26606 38113
rect 26290 38048 26296 38112
rect 26360 38048 26376 38112
rect 26440 38048 26456 38112
rect 26520 38048 26536 38112
rect 26600 38048 26606 38112
rect 26290 38047 26606 38048
rect 35200 38028 36000 38118
rect 0 37498 800 37588
rect 5170 37568 5486 37569
rect 5170 37504 5176 37568
rect 5240 37504 5256 37568
rect 5320 37504 5336 37568
rect 5400 37504 5416 37568
rect 5480 37504 5486 37568
rect 5170 37503 5486 37504
rect 13618 37568 13934 37569
rect 13618 37504 13624 37568
rect 13688 37504 13704 37568
rect 13768 37504 13784 37568
rect 13848 37504 13864 37568
rect 13928 37504 13934 37568
rect 13618 37503 13934 37504
rect 22066 37568 22382 37569
rect 22066 37504 22072 37568
rect 22136 37504 22152 37568
rect 22216 37504 22232 37568
rect 22296 37504 22312 37568
rect 22376 37504 22382 37568
rect 22066 37503 22382 37504
rect 30514 37568 30830 37569
rect 30514 37504 30520 37568
rect 30584 37504 30600 37568
rect 30664 37504 30680 37568
rect 30744 37504 30760 37568
rect 30824 37504 30830 37568
rect 30514 37503 30830 37504
rect 3325 37498 3391 37501
rect 0 37496 3391 37498
rect 0 37440 3330 37496
rect 3386 37440 3391 37496
rect 0 37438 3391 37440
rect 0 37348 800 37438
rect 3325 37435 3391 37438
rect 35200 37348 36000 37588
rect 9394 37024 9710 37025
rect 9394 36960 9400 37024
rect 9464 36960 9480 37024
rect 9544 36960 9560 37024
rect 9624 36960 9640 37024
rect 9704 36960 9710 37024
rect 9394 36959 9710 36960
rect 17842 37024 18158 37025
rect 17842 36960 17848 37024
rect 17912 36960 17928 37024
rect 17992 36960 18008 37024
rect 18072 36960 18088 37024
rect 18152 36960 18158 37024
rect 17842 36959 18158 36960
rect 26290 37024 26606 37025
rect 26290 36960 26296 37024
rect 26360 36960 26376 37024
rect 26440 36960 26456 37024
rect 26520 36960 26536 37024
rect 26600 36960 26606 37024
rect 26290 36959 26606 36960
rect 0 36818 800 36908
rect 4061 36818 4127 36821
rect 0 36816 4127 36818
rect 0 36760 4066 36816
rect 4122 36760 4127 36816
rect 0 36758 4127 36760
rect 0 36668 800 36758
rect 4061 36755 4127 36758
rect 31661 36818 31727 36821
rect 35200 36818 36000 36908
rect 31661 36816 36000 36818
rect 31661 36760 31666 36816
rect 31722 36760 36000 36816
rect 31661 36758 36000 36760
rect 31661 36755 31727 36758
rect 35200 36668 36000 36758
rect 5170 36480 5486 36481
rect 5170 36416 5176 36480
rect 5240 36416 5256 36480
rect 5320 36416 5336 36480
rect 5400 36416 5416 36480
rect 5480 36416 5486 36480
rect 5170 36415 5486 36416
rect 13618 36480 13934 36481
rect 13618 36416 13624 36480
rect 13688 36416 13704 36480
rect 13768 36416 13784 36480
rect 13848 36416 13864 36480
rect 13928 36416 13934 36480
rect 13618 36415 13934 36416
rect 22066 36480 22382 36481
rect 22066 36416 22072 36480
rect 22136 36416 22152 36480
rect 22216 36416 22232 36480
rect 22296 36416 22312 36480
rect 22376 36416 22382 36480
rect 22066 36415 22382 36416
rect 30514 36480 30830 36481
rect 30514 36416 30520 36480
rect 30584 36416 30600 36480
rect 30664 36416 30680 36480
rect 30744 36416 30760 36480
rect 30824 36416 30830 36480
rect 30514 36415 30830 36416
rect 0 36138 800 36228
rect 1853 36138 1919 36141
rect 0 36136 1919 36138
rect 0 36080 1858 36136
rect 1914 36080 1919 36136
rect 0 36078 1919 36080
rect 0 35988 800 36078
rect 1853 36075 1919 36078
rect 35200 35988 36000 36228
rect 9394 35936 9710 35937
rect 9394 35872 9400 35936
rect 9464 35872 9480 35936
rect 9544 35872 9560 35936
rect 9624 35872 9640 35936
rect 9704 35872 9710 35936
rect 9394 35871 9710 35872
rect 17842 35936 18158 35937
rect 17842 35872 17848 35936
rect 17912 35872 17928 35936
rect 17992 35872 18008 35936
rect 18072 35872 18088 35936
rect 18152 35872 18158 35936
rect 17842 35871 18158 35872
rect 26290 35936 26606 35937
rect 26290 35872 26296 35936
rect 26360 35872 26376 35936
rect 26440 35872 26456 35936
rect 26520 35872 26536 35936
rect 26600 35872 26606 35936
rect 26290 35871 26606 35872
rect 0 35458 800 35548
rect 3325 35458 3391 35461
rect 0 35456 3391 35458
rect 0 35400 3330 35456
rect 3386 35400 3391 35456
rect 0 35398 3391 35400
rect 0 35308 800 35398
rect 3325 35395 3391 35398
rect 5170 35392 5486 35393
rect 5170 35328 5176 35392
rect 5240 35328 5256 35392
rect 5320 35328 5336 35392
rect 5400 35328 5416 35392
rect 5480 35328 5486 35392
rect 5170 35327 5486 35328
rect 13618 35392 13934 35393
rect 13618 35328 13624 35392
rect 13688 35328 13704 35392
rect 13768 35328 13784 35392
rect 13848 35328 13864 35392
rect 13928 35328 13934 35392
rect 13618 35327 13934 35328
rect 22066 35392 22382 35393
rect 22066 35328 22072 35392
rect 22136 35328 22152 35392
rect 22216 35328 22232 35392
rect 22296 35328 22312 35392
rect 22376 35328 22382 35392
rect 22066 35327 22382 35328
rect 30514 35392 30830 35393
rect 30514 35328 30520 35392
rect 30584 35328 30600 35392
rect 30664 35328 30680 35392
rect 30744 35328 30760 35392
rect 30824 35328 30830 35392
rect 30514 35327 30830 35328
rect 0 34628 800 34868
rect 9394 34848 9710 34849
rect 9394 34784 9400 34848
rect 9464 34784 9480 34848
rect 9544 34784 9560 34848
rect 9624 34784 9640 34848
rect 9704 34784 9710 34848
rect 9394 34783 9710 34784
rect 17842 34848 18158 34849
rect 17842 34784 17848 34848
rect 17912 34784 17928 34848
rect 17992 34784 18008 34848
rect 18072 34784 18088 34848
rect 18152 34784 18158 34848
rect 17842 34783 18158 34784
rect 26290 34848 26606 34849
rect 26290 34784 26296 34848
rect 26360 34784 26376 34848
rect 26440 34784 26456 34848
rect 26520 34784 26536 34848
rect 26600 34784 26606 34848
rect 26290 34783 26606 34784
rect 31569 34778 31635 34781
rect 35200 34778 36000 34868
rect 31569 34776 36000 34778
rect 31569 34720 31574 34776
rect 31630 34720 36000 34776
rect 31569 34718 36000 34720
rect 31569 34715 31635 34718
rect 35200 34628 36000 34718
rect 5170 34304 5486 34305
rect 5170 34240 5176 34304
rect 5240 34240 5256 34304
rect 5320 34240 5336 34304
rect 5400 34240 5416 34304
rect 5480 34240 5486 34304
rect 5170 34239 5486 34240
rect 13618 34304 13934 34305
rect 13618 34240 13624 34304
rect 13688 34240 13704 34304
rect 13768 34240 13784 34304
rect 13848 34240 13864 34304
rect 13928 34240 13934 34304
rect 13618 34239 13934 34240
rect 22066 34304 22382 34305
rect 22066 34240 22072 34304
rect 22136 34240 22152 34304
rect 22216 34240 22232 34304
rect 22296 34240 22312 34304
rect 22376 34240 22382 34304
rect 22066 34239 22382 34240
rect 30514 34304 30830 34305
rect 30514 34240 30520 34304
rect 30584 34240 30600 34304
rect 30664 34240 30680 34304
rect 30744 34240 30760 34304
rect 30824 34240 30830 34304
rect 30514 34239 30830 34240
rect 0 34098 800 34188
rect 3417 34098 3483 34101
rect 0 34096 3483 34098
rect 0 34040 3422 34096
rect 3478 34040 3483 34096
rect 0 34038 3483 34040
rect 0 33948 800 34038
rect 3417 34035 3483 34038
rect 32949 34098 33015 34101
rect 35200 34098 36000 34188
rect 32949 34096 36000 34098
rect 32949 34040 32954 34096
rect 33010 34040 36000 34096
rect 32949 34038 36000 34040
rect 32949 34035 33015 34038
rect 35200 33948 36000 34038
rect 9394 33760 9710 33761
rect 9394 33696 9400 33760
rect 9464 33696 9480 33760
rect 9544 33696 9560 33760
rect 9624 33696 9640 33760
rect 9704 33696 9710 33760
rect 9394 33695 9710 33696
rect 17842 33760 18158 33761
rect 17842 33696 17848 33760
rect 17912 33696 17928 33760
rect 17992 33696 18008 33760
rect 18072 33696 18088 33760
rect 18152 33696 18158 33760
rect 17842 33695 18158 33696
rect 26290 33760 26606 33761
rect 26290 33696 26296 33760
rect 26360 33696 26376 33760
rect 26440 33696 26456 33760
rect 26520 33696 26536 33760
rect 26600 33696 26606 33760
rect 26290 33695 26606 33696
rect 32305 33418 32371 33421
rect 35200 33418 36000 33508
rect 32305 33416 36000 33418
rect 32305 33360 32310 33416
rect 32366 33360 36000 33416
rect 32305 33358 36000 33360
rect 32305 33355 32371 33358
rect 35200 33268 36000 33358
rect 5170 33216 5486 33217
rect 5170 33152 5176 33216
rect 5240 33152 5256 33216
rect 5320 33152 5336 33216
rect 5400 33152 5416 33216
rect 5480 33152 5486 33216
rect 5170 33151 5486 33152
rect 13618 33216 13934 33217
rect 13618 33152 13624 33216
rect 13688 33152 13704 33216
rect 13768 33152 13784 33216
rect 13848 33152 13864 33216
rect 13928 33152 13934 33216
rect 13618 33151 13934 33152
rect 22066 33216 22382 33217
rect 22066 33152 22072 33216
rect 22136 33152 22152 33216
rect 22216 33152 22232 33216
rect 22296 33152 22312 33216
rect 22376 33152 22382 33216
rect 22066 33151 22382 33152
rect 30514 33216 30830 33217
rect 30514 33152 30520 33216
rect 30584 33152 30600 33216
rect 30664 33152 30680 33216
rect 30744 33152 30760 33216
rect 30824 33152 30830 33216
rect 30514 33151 30830 33152
rect 0 32588 800 32828
rect 33685 32738 33751 32741
rect 35200 32738 36000 32828
rect 33685 32736 36000 32738
rect 33685 32680 33690 32736
rect 33746 32680 36000 32736
rect 33685 32678 36000 32680
rect 33685 32675 33751 32678
rect 9394 32672 9710 32673
rect 9394 32608 9400 32672
rect 9464 32608 9480 32672
rect 9544 32608 9560 32672
rect 9624 32608 9640 32672
rect 9704 32608 9710 32672
rect 9394 32607 9710 32608
rect 17842 32672 18158 32673
rect 17842 32608 17848 32672
rect 17912 32608 17928 32672
rect 17992 32608 18008 32672
rect 18072 32608 18088 32672
rect 18152 32608 18158 32672
rect 17842 32607 18158 32608
rect 26290 32672 26606 32673
rect 26290 32608 26296 32672
rect 26360 32608 26376 32672
rect 26440 32608 26456 32672
rect 26520 32608 26536 32672
rect 26600 32608 26606 32672
rect 26290 32607 26606 32608
rect 35200 32588 36000 32678
rect 0 32058 800 32148
rect 5170 32128 5486 32129
rect 5170 32064 5176 32128
rect 5240 32064 5256 32128
rect 5320 32064 5336 32128
rect 5400 32064 5416 32128
rect 5480 32064 5486 32128
rect 5170 32063 5486 32064
rect 13618 32128 13934 32129
rect 13618 32064 13624 32128
rect 13688 32064 13704 32128
rect 13768 32064 13784 32128
rect 13848 32064 13864 32128
rect 13928 32064 13934 32128
rect 13618 32063 13934 32064
rect 22066 32128 22382 32129
rect 22066 32064 22072 32128
rect 22136 32064 22152 32128
rect 22216 32064 22232 32128
rect 22296 32064 22312 32128
rect 22376 32064 22382 32128
rect 22066 32063 22382 32064
rect 30514 32128 30830 32129
rect 30514 32064 30520 32128
rect 30584 32064 30600 32128
rect 30664 32064 30680 32128
rect 30744 32064 30760 32128
rect 30824 32064 30830 32128
rect 30514 32063 30830 32064
rect 3417 32058 3483 32061
rect 0 32056 3483 32058
rect 0 32000 3422 32056
rect 3478 32000 3483 32056
rect 0 31998 3483 32000
rect 0 31908 800 31998
rect 3417 31995 3483 31998
rect 33041 32058 33107 32061
rect 35200 32058 36000 32148
rect 33041 32056 36000 32058
rect 33041 32000 33046 32056
rect 33102 32000 36000 32056
rect 33041 31998 36000 32000
rect 33041 31995 33107 31998
rect 35200 31908 36000 31998
rect 9394 31584 9710 31585
rect 9394 31520 9400 31584
rect 9464 31520 9480 31584
rect 9544 31520 9560 31584
rect 9624 31520 9640 31584
rect 9704 31520 9710 31584
rect 9394 31519 9710 31520
rect 17842 31584 18158 31585
rect 17842 31520 17848 31584
rect 17912 31520 17928 31584
rect 17992 31520 18008 31584
rect 18072 31520 18088 31584
rect 18152 31520 18158 31584
rect 17842 31519 18158 31520
rect 26290 31584 26606 31585
rect 26290 31520 26296 31584
rect 26360 31520 26376 31584
rect 26440 31520 26456 31584
rect 26520 31520 26536 31584
rect 26600 31520 26606 31584
rect 26290 31519 26606 31520
rect 0 31378 800 31468
rect 3417 31378 3483 31381
rect 0 31376 3483 31378
rect 0 31320 3422 31376
rect 3478 31320 3483 31376
rect 0 31318 3483 31320
rect 0 31228 800 31318
rect 3417 31315 3483 31318
rect 34145 31378 34211 31381
rect 35200 31378 36000 31468
rect 34145 31376 36000 31378
rect 34145 31320 34150 31376
rect 34206 31320 36000 31376
rect 34145 31318 36000 31320
rect 34145 31315 34211 31318
rect 35200 31228 36000 31318
rect 5170 31040 5486 31041
rect 5170 30976 5176 31040
rect 5240 30976 5256 31040
rect 5320 30976 5336 31040
rect 5400 30976 5416 31040
rect 5480 30976 5486 31040
rect 5170 30975 5486 30976
rect 13618 31040 13934 31041
rect 13618 30976 13624 31040
rect 13688 30976 13704 31040
rect 13768 30976 13784 31040
rect 13848 30976 13864 31040
rect 13928 30976 13934 31040
rect 13618 30975 13934 30976
rect 22066 31040 22382 31041
rect 22066 30976 22072 31040
rect 22136 30976 22152 31040
rect 22216 30976 22232 31040
rect 22296 30976 22312 31040
rect 22376 30976 22382 31040
rect 22066 30975 22382 30976
rect 30514 31040 30830 31041
rect 30514 30976 30520 31040
rect 30584 30976 30600 31040
rect 30664 30976 30680 31040
rect 30744 30976 30760 31040
rect 30824 30976 30830 31040
rect 30514 30975 30830 30976
rect 0 30548 800 30788
rect 35200 30548 36000 30788
rect 9394 30496 9710 30497
rect 9394 30432 9400 30496
rect 9464 30432 9480 30496
rect 9544 30432 9560 30496
rect 9624 30432 9640 30496
rect 9704 30432 9710 30496
rect 9394 30431 9710 30432
rect 17842 30496 18158 30497
rect 17842 30432 17848 30496
rect 17912 30432 17928 30496
rect 17992 30432 18008 30496
rect 18072 30432 18088 30496
rect 18152 30432 18158 30496
rect 17842 30431 18158 30432
rect 26290 30496 26606 30497
rect 26290 30432 26296 30496
rect 26360 30432 26376 30496
rect 26440 30432 26456 30496
rect 26520 30432 26536 30496
rect 26600 30432 26606 30496
rect 26290 30431 26606 30432
rect 0 29868 800 30108
rect 5170 29952 5486 29953
rect 5170 29888 5176 29952
rect 5240 29888 5256 29952
rect 5320 29888 5336 29952
rect 5400 29888 5416 29952
rect 5480 29888 5486 29952
rect 5170 29887 5486 29888
rect 13618 29952 13934 29953
rect 13618 29888 13624 29952
rect 13688 29888 13704 29952
rect 13768 29888 13784 29952
rect 13848 29888 13864 29952
rect 13928 29888 13934 29952
rect 13618 29887 13934 29888
rect 22066 29952 22382 29953
rect 22066 29888 22072 29952
rect 22136 29888 22152 29952
rect 22216 29888 22232 29952
rect 22296 29888 22312 29952
rect 22376 29888 22382 29952
rect 22066 29887 22382 29888
rect 30514 29952 30830 29953
rect 30514 29888 30520 29952
rect 30584 29888 30600 29952
rect 30664 29888 30680 29952
rect 30744 29888 30760 29952
rect 30824 29888 30830 29952
rect 30514 29887 30830 29888
rect 35200 29868 36000 30108
rect 0 29188 800 29428
rect 9394 29408 9710 29409
rect 9394 29344 9400 29408
rect 9464 29344 9480 29408
rect 9544 29344 9560 29408
rect 9624 29344 9640 29408
rect 9704 29344 9710 29408
rect 9394 29343 9710 29344
rect 17842 29408 18158 29409
rect 17842 29344 17848 29408
rect 17912 29344 17928 29408
rect 17992 29344 18008 29408
rect 18072 29344 18088 29408
rect 18152 29344 18158 29408
rect 17842 29343 18158 29344
rect 26290 29408 26606 29409
rect 26290 29344 26296 29408
rect 26360 29344 26376 29408
rect 26440 29344 26456 29408
rect 26520 29344 26536 29408
rect 26600 29344 26606 29408
rect 26290 29343 26606 29344
rect 35200 29188 36000 29428
rect 5170 28864 5486 28865
rect 5170 28800 5176 28864
rect 5240 28800 5256 28864
rect 5320 28800 5336 28864
rect 5400 28800 5416 28864
rect 5480 28800 5486 28864
rect 5170 28799 5486 28800
rect 13618 28864 13934 28865
rect 13618 28800 13624 28864
rect 13688 28800 13704 28864
rect 13768 28800 13784 28864
rect 13848 28800 13864 28864
rect 13928 28800 13934 28864
rect 13618 28799 13934 28800
rect 22066 28864 22382 28865
rect 22066 28800 22072 28864
rect 22136 28800 22152 28864
rect 22216 28800 22232 28864
rect 22296 28800 22312 28864
rect 22376 28800 22382 28864
rect 22066 28799 22382 28800
rect 30514 28864 30830 28865
rect 30514 28800 30520 28864
rect 30584 28800 30600 28864
rect 30664 28800 30680 28864
rect 30744 28800 30760 28864
rect 30824 28800 30830 28864
rect 30514 28799 30830 28800
rect 0 28508 800 28748
rect 9394 28320 9710 28321
rect 9394 28256 9400 28320
rect 9464 28256 9480 28320
rect 9544 28256 9560 28320
rect 9624 28256 9640 28320
rect 9704 28256 9710 28320
rect 9394 28255 9710 28256
rect 17842 28320 18158 28321
rect 17842 28256 17848 28320
rect 17912 28256 17928 28320
rect 17992 28256 18008 28320
rect 18072 28256 18088 28320
rect 18152 28256 18158 28320
rect 17842 28255 18158 28256
rect 26290 28320 26606 28321
rect 26290 28256 26296 28320
rect 26360 28256 26376 28320
rect 26440 28256 26456 28320
rect 26520 28256 26536 28320
rect 26600 28256 26606 28320
rect 26290 28255 26606 28256
rect 0 27828 800 28068
rect 33041 27978 33107 27981
rect 35200 27978 36000 28068
rect 33041 27976 36000 27978
rect 33041 27920 33046 27976
rect 33102 27920 36000 27976
rect 33041 27918 36000 27920
rect 33041 27915 33107 27918
rect 35200 27828 36000 27918
rect 5170 27776 5486 27777
rect 5170 27712 5176 27776
rect 5240 27712 5256 27776
rect 5320 27712 5336 27776
rect 5400 27712 5416 27776
rect 5480 27712 5486 27776
rect 5170 27711 5486 27712
rect 13618 27776 13934 27777
rect 13618 27712 13624 27776
rect 13688 27712 13704 27776
rect 13768 27712 13784 27776
rect 13848 27712 13864 27776
rect 13928 27712 13934 27776
rect 13618 27711 13934 27712
rect 22066 27776 22382 27777
rect 22066 27712 22072 27776
rect 22136 27712 22152 27776
rect 22216 27712 22232 27776
rect 22296 27712 22312 27776
rect 22376 27712 22382 27776
rect 22066 27711 22382 27712
rect 30514 27776 30830 27777
rect 30514 27712 30520 27776
rect 30584 27712 30600 27776
rect 30664 27712 30680 27776
rect 30744 27712 30760 27776
rect 30824 27712 30830 27776
rect 30514 27711 30830 27712
rect 0 27148 800 27388
rect 9394 27232 9710 27233
rect 9394 27168 9400 27232
rect 9464 27168 9480 27232
rect 9544 27168 9560 27232
rect 9624 27168 9640 27232
rect 9704 27168 9710 27232
rect 9394 27167 9710 27168
rect 17842 27232 18158 27233
rect 17842 27168 17848 27232
rect 17912 27168 17928 27232
rect 17992 27168 18008 27232
rect 18072 27168 18088 27232
rect 18152 27168 18158 27232
rect 17842 27167 18158 27168
rect 26290 27232 26606 27233
rect 26290 27168 26296 27232
rect 26360 27168 26376 27232
rect 26440 27168 26456 27232
rect 26520 27168 26536 27232
rect 26600 27168 26606 27232
rect 26290 27167 26606 27168
rect 35200 27148 36000 27388
rect 5170 26688 5486 26689
rect 5170 26624 5176 26688
rect 5240 26624 5256 26688
rect 5320 26624 5336 26688
rect 5400 26624 5416 26688
rect 5480 26624 5486 26688
rect 5170 26623 5486 26624
rect 13618 26688 13934 26689
rect 13618 26624 13624 26688
rect 13688 26624 13704 26688
rect 13768 26624 13784 26688
rect 13848 26624 13864 26688
rect 13928 26624 13934 26688
rect 13618 26623 13934 26624
rect 22066 26688 22382 26689
rect 22066 26624 22072 26688
rect 22136 26624 22152 26688
rect 22216 26624 22232 26688
rect 22296 26624 22312 26688
rect 22376 26624 22382 26688
rect 22066 26623 22382 26624
rect 30514 26688 30830 26689
rect 30514 26624 30520 26688
rect 30584 26624 30600 26688
rect 30664 26624 30680 26688
rect 30744 26624 30760 26688
rect 30824 26624 30830 26688
rect 30514 26623 30830 26624
rect 35200 26468 36000 26708
rect 9394 26144 9710 26145
rect 9394 26080 9400 26144
rect 9464 26080 9480 26144
rect 9544 26080 9560 26144
rect 9624 26080 9640 26144
rect 9704 26080 9710 26144
rect 9394 26079 9710 26080
rect 17842 26144 18158 26145
rect 17842 26080 17848 26144
rect 17912 26080 17928 26144
rect 17992 26080 18008 26144
rect 18072 26080 18088 26144
rect 18152 26080 18158 26144
rect 17842 26079 18158 26080
rect 26290 26144 26606 26145
rect 26290 26080 26296 26144
rect 26360 26080 26376 26144
rect 26440 26080 26456 26144
rect 26520 26080 26536 26144
rect 26600 26080 26606 26144
rect 26290 26079 26606 26080
rect 0 25788 800 26028
rect 33041 25938 33107 25941
rect 35200 25938 36000 26028
rect 33041 25936 36000 25938
rect 33041 25880 33046 25936
rect 33102 25880 36000 25936
rect 33041 25878 36000 25880
rect 33041 25875 33107 25878
rect 35200 25788 36000 25878
rect 5170 25600 5486 25601
rect 5170 25536 5176 25600
rect 5240 25536 5256 25600
rect 5320 25536 5336 25600
rect 5400 25536 5416 25600
rect 5480 25536 5486 25600
rect 5170 25535 5486 25536
rect 13618 25600 13934 25601
rect 13618 25536 13624 25600
rect 13688 25536 13704 25600
rect 13768 25536 13784 25600
rect 13848 25536 13864 25600
rect 13928 25536 13934 25600
rect 13618 25535 13934 25536
rect 22066 25600 22382 25601
rect 22066 25536 22072 25600
rect 22136 25536 22152 25600
rect 22216 25536 22232 25600
rect 22296 25536 22312 25600
rect 22376 25536 22382 25600
rect 22066 25535 22382 25536
rect 30514 25600 30830 25601
rect 30514 25536 30520 25600
rect 30584 25536 30600 25600
rect 30664 25536 30680 25600
rect 30744 25536 30760 25600
rect 30824 25536 30830 25600
rect 30514 25535 30830 25536
rect 0 25258 800 25348
rect 3417 25258 3483 25261
rect 0 25256 3483 25258
rect 0 25200 3422 25256
rect 3478 25200 3483 25256
rect 0 25198 3483 25200
rect 0 25108 800 25198
rect 3417 25195 3483 25198
rect 31753 25258 31819 25261
rect 35200 25258 36000 25348
rect 31753 25256 36000 25258
rect 31753 25200 31758 25256
rect 31814 25200 36000 25256
rect 31753 25198 36000 25200
rect 31753 25195 31819 25198
rect 35200 25108 36000 25198
rect 9394 25056 9710 25057
rect 9394 24992 9400 25056
rect 9464 24992 9480 25056
rect 9544 24992 9560 25056
rect 9624 24992 9640 25056
rect 9704 24992 9710 25056
rect 9394 24991 9710 24992
rect 17842 25056 18158 25057
rect 17842 24992 17848 25056
rect 17912 24992 17928 25056
rect 17992 24992 18008 25056
rect 18072 24992 18088 25056
rect 18152 24992 18158 25056
rect 17842 24991 18158 24992
rect 26290 25056 26606 25057
rect 26290 24992 26296 25056
rect 26360 24992 26376 25056
rect 26440 24992 26456 25056
rect 26520 24992 26536 25056
rect 26600 24992 26606 25056
rect 26290 24991 26606 24992
rect 0 24428 800 24668
rect 32673 24578 32739 24581
rect 35200 24578 36000 24668
rect 32673 24576 36000 24578
rect 32673 24520 32678 24576
rect 32734 24520 36000 24576
rect 32673 24518 36000 24520
rect 32673 24515 32739 24518
rect 5170 24512 5486 24513
rect 5170 24448 5176 24512
rect 5240 24448 5256 24512
rect 5320 24448 5336 24512
rect 5400 24448 5416 24512
rect 5480 24448 5486 24512
rect 5170 24447 5486 24448
rect 13618 24512 13934 24513
rect 13618 24448 13624 24512
rect 13688 24448 13704 24512
rect 13768 24448 13784 24512
rect 13848 24448 13864 24512
rect 13928 24448 13934 24512
rect 13618 24447 13934 24448
rect 22066 24512 22382 24513
rect 22066 24448 22072 24512
rect 22136 24448 22152 24512
rect 22216 24448 22232 24512
rect 22296 24448 22312 24512
rect 22376 24448 22382 24512
rect 22066 24447 22382 24448
rect 30514 24512 30830 24513
rect 30514 24448 30520 24512
rect 30584 24448 30600 24512
rect 30664 24448 30680 24512
rect 30744 24448 30760 24512
rect 30824 24448 30830 24512
rect 30514 24447 30830 24448
rect 35200 24428 36000 24518
rect 0 23748 800 23988
rect 9394 23968 9710 23969
rect 9394 23904 9400 23968
rect 9464 23904 9480 23968
rect 9544 23904 9560 23968
rect 9624 23904 9640 23968
rect 9704 23904 9710 23968
rect 9394 23903 9710 23904
rect 17842 23968 18158 23969
rect 17842 23904 17848 23968
rect 17912 23904 17928 23968
rect 17992 23904 18008 23968
rect 18072 23904 18088 23968
rect 18152 23904 18158 23968
rect 17842 23903 18158 23904
rect 26290 23968 26606 23969
rect 26290 23904 26296 23968
rect 26360 23904 26376 23968
rect 26440 23904 26456 23968
rect 26520 23904 26536 23968
rect 26600 23904 26606 23968
rect 26290 23903 26606 23904
rect 34145 23898 34211 23901
rect 35200 23898 36000 23988
rect 34145 23896 36000 23898
rect 34145 23840 34150 23896
rect 34206 23840 36000 23896
rect 34145 23838 36000 23840
rect 34145 23835 34211 23838
rect 35200 23748 36000 23838
rect 5170 23424 5486 23425
rect 5170 23360 5176 23424
rect 5240 23360 5256 23424
rect 5320 23360 5336 23424
rect 5400 23360 5416 23424
rect 5480 23360 5486 23424
rect 5170 23359 5486 23360
rect 13618 23424 13934 23425
rect 13618 23360 13624 23424
rect 13688 23360 13704 23424
rect 13768 23360 13784 23424
rect 13848 23360 13864 23424
rect 13928 23360 13934 23424
rect 13618 23359 13934 23360
rect 22066 23424 22382 23425
rect 22066 23360 22072 23424
rect 22136 23360 22152 23424
rect 22216 23360 22232 23424
rect 22296 23360 22312 23424
rect 22376 23360 22382 23424
rect 22066 23359 22382 23360
rect 30514 23424 30830 23425
rect 30514 23360 30520 23424
rect 30584 23360 30600 23424
rect 30664 23360 30680 23424
rect 30744 23360 30760 23424
rect 30824 23360 30830 23424
rect 30514 23359 30830 23360
rect 0 23068 800 23308
rect 34145 23218 34211 23221
rect 35200 23218 36000 23308
rect 34145 23216 36000 23218
rect 34145 23160 34150 23216
rect 34206 23160 36000 23216
rect 34145 23158 36000 23160
rect 34145 23155 34211 23158
rect 35200 23068 36000 23158
rect 9394 22880 9710 22881
rect 9394 22816 9400 22880
rect 9464 22816 9480 22880
rect 9544 22816 9560 22880
rect 9624 22816 9640 22880
rect 9704 22816 9710 22880
rect 9394 22815 9710 22816
rect 17842 22880 18158 22881
rect 17842 22816 17848 22880
rect 17912 22816 17928 22880
rect 17992 22816 18008 22880
rect 18072 22816 18088 22880
rect 18152 22816 18158 22880
rect 17842 22815 18158 22816
rect 26290 22880 26606 22881
rect 26290 22816 26296 22880
rect 26360 22816 26376 22880
rect 26440 22816 26456 22880
rect 26520 22816 26536 22880
rect 26600 22816 26606 22880
rect 26290 22815 26606 22816
rect 0 22388 800 22628
rect 35200 22388 36000 22628
rect 5170 22336 5486 22337
rect 5170 22272 5176 22336
rect 5240 22272 5256 22336
rect 5320 22272 5336 22336
rect 5400 22272 5416 22336
rect 5480 22272 5486 22336
rect 5170 22271 5486 22272
rect 13618 22336 13934 22337
rect 13618 22272 13624 22336
rect 13688 22272 13704 22336
rect 13768 22272 13784 22336
rect 13848 22272 13864 22336
rect 13928 22272 13934 22336
rect 13618 22271 13934 22272
rect 22066 22336 22382 22337
rect 22066 22272 22072 22336
rect 22136 22272 22152 22336
rect 22216 22272 22232 22336
rect 22296 22272 22312 22336
rect 22376 22272 22382 22336
rect 22066 22271 22382 22272
rect 30514 22336 30830 22337
rect 30514 22272 30520 22336
rect 30584 22272 30600 22336
rect 30664 22272 30680 22336
rect 30744 22272 30760 22336
rect 30824 22272 30830 22336
rect 30514 22271 30830 22272
rect 0 21708 800 21948
rect 9394 21792 9710 21793
rect 9394 21728 9400 21792
rect 9464 21728 9480 21792
rect 9544 21728 9560 21792
rect 9624 21728 9640 21792
rect 9704 21728 9710 21792
rect 9394 21727 9710 21728
rect 17842 21792 18158 21793
rect 17842 21728 17848 21792
rect 17912 21728 17928 21792
rect 17992 21728 18008 21792
rect 18072 21728 18088 21792
rect 18152 21728 18158 21792
rect 17842 21727 18158 21728
rect 26290 21792 26606 21793
rect 26290 21728 26296 21792
rect 26360 21728 26376 21792
rect 26440 21728 26456 21792
rect 26520 21728 26536 21792
rect 26600 21728 26606 21792
rect 26290 21727 26606 21728
rect 0 21028 800 21268
rect 5170 21248 5486 21249
rect 5170 21184 5176 21248
rect 5240 21184 5256 21248
rect 5320 21184 5336 21248
rect 5400 21184 5416 21248
rect 5480 21184 5486 21248
rect 5170 21183 5486 21184
rect 13618 21248 13934 21249
rect 13618 21184 13624 21248
rect 13688 21184 13704 21248
rect 13768 21184 13784 21248
rect 13848 21184 13864 21248
rect 13928 21184 13934 21248
rect 13618 21183 13934 21184
rect 22066 21248 22382 21249
rect 22066 21184 22072 21248
rect 22136 21184 22152 21248
rect 22216 21184 22232 21248
rect 22296 21184 22312 21248
rect 22376 21184 22382 21248
rect 22066 21183 22382 21184
rect 30514 21248 30830 21249
rect 30514 21184 30520 21248
rect 30584 21184 30600 21248
rect 30664 21184 30680 21248
rect 30744 21184 30760 21248
rect 30824 21184 30830 21248
rect 30514 21183 30830 21184
rect 35200 21028 36000 21268
rect 9394 20704 9710 20705
rect 9394 20640 9400 20704
rect 9464 20640 9480 20704
rect 9544 20640 9560 20704
rect 9624 20640 9640 20704
rect 9704 20640 9710 20704
rect 9394 20639 9710 20640
rect 17842 20704 18158 20705
rect 17842 20640 17848 20704
rect 17912 20640 17928 20704
rect 17992 20640 18008 20704
rect 18072 20640 18088 20704
rect 18152 20640 18158 20704
rect 17842 20639 18158 20640
rect 26290 20704 26606 20705
rect 26290 20640 26296 20704
rect 26360 20640 26376 20704
rect 26440 20640 26456 20704
rect 26520 20640 26536 20704
rect 26600 20640 26606 20704
rect 26290 20639 26606 20640
rect 0 20348 800 20588
rect 32949 20498 33015 20501
rect 35200 20498 36000 20588
rect 32949 20496 36000 20498
rect 32949 20440 32954 20496
rect 33010 20440 36000 20496
rect 32949 20438 36000 20440
rect 32949 20435 33015 20438
rect 35200 20348 36000 20438
rect 5170 20160 5486 20161
rect 5170 20096 5176 20160
rect 5240 20096 5256 20160
rect 5320 20096 5336 20160
rect 5400 20096 5416 20160
rect 5480 20096 5486 20160
rect 5170 20095 5486 20096
rect 13618 20160 13934 20161
rect 13618 20096 13624 20160
rect 13688 20096 13704 20160
rect 13768 20096 13784 20160
rect 13848 20096 13864 20160
rect 13928 20096 13934 20160
rect 13618 20095 13934 20096
rect 22066 20160 22382 20161
rect 22066 20096 22072 20160
rect 22136 20096 22152 20160
rect 22216 20096 22232 20160
rect 22296 20096 22312 20160
rect 22376 20096 22382 20160
rect 22066 20095 22382 20096
rect 30514 20160 30830 20161
rect 30514 20096 30520 20160
rect 30584 20096 30600 20160
rect 30664 20096 30680 20160
rect 30744 20096 30760 20160
rect 30824 20096 30830 20160
rect 30514 20095 30830 20096
rect 31753 19818 31819 19821
rect 35200 19818 36000 19908
rect 31753 19816 36000 19818
rect 31753 19760 31758 19816
rect 31814 19760 36000 19816
rect 31753 19758 36000 19760
rect 31753 19755 31819 19758
rect 35200 19668 36000 19758
rect 9394 19616 9710 19617
rect 9394 19552 9400 19616
rect 9464 19552 9480 19616
rect 9544 19552 9560 19616
rect 9624 19552 9640 19616
rect 9704 19552 9710 19616
rect 9394 19551 9710 19552
rect 17842 19616 18158 19617
rect 17842 19552 17848 19616
rect 17912 19552 17928 19616
rect 17992 19552 18008 19616
rect 18072 19552 18088 19616
rect 18152 19552 18158 19616
rect 17842 19551 18158 19552
rect 26290 19616 26606 19617
rect 26290 19552 26296 19616
rect 26360 19552 26376 19616
rect 26440 19552 26456 19616
rect 26520 19552 26536 19616
rect 26600 19552 26606 19616
rect 26290 19551 26606 19552
rect 0 19138 800 19228
rect 3417 19138 3483 19141
rect 0 19136 3483 19138
rect 0 19080 3422 19136
rect 3478 19080 3483 19136
rect 0 19078 3483 19080
rect 0 18988 800 19078
rect 3417 19075 3483 19078
rect 33041 19138 33107 19141
rect 35200 19138 36000 19228
rect 33041 19136 36000 19138
rect 33041 19080 33046 19136
rect 33102 19080 36000 19136
rect 33041 19078 36000 19080
rect 33041 19075 33107 19078
rect 5170 19072 5486 19073
rect 5170 19008 5176 19072
rect 5240 19008 5256 19072
rect 5320 19008 5336 19072
rect 5400 19008 5416 19072
rect 5480 19008 5486 19072
rect 5170 19007 5486 19008
rect 13618 19072 13934 19073
rect 13618 19008 13624 19072
rect 13688 19008 13704 19072
rect 13768 19008 13784 19072
rect 13848 19008 13864 19072
rect 13928 19008 13934 19072
rect 13618 19007 13934 19008
rect 22066 19072 22382 19073
rect 22066 19008 22072 19072
rect 22136 19008 22152 19072
rect 22216 19008 22232 19072
rect 22296 19008 22312 19072
rect 22376 19008 22382 19072
rect 22066 19007 22382 19008
rect 30514 19072 30830 19073
rect 30514 19008 30520 19072
rect 30584 19008 30600 19072
rect 30664 19008 30680 19072
rect 30744 19008 30760 19072
rect 30824 19008 30830 19072
rect 30514 19007 30830 19008
rect 35200 18988 36000 19078
rect 0 18458 800 18548
rect 9394 18528 9710 18529
rect 9394 18464 9400 18528
rect 9464 18464 9480 18528
rect 9544 18464 9560 18528
rect 9624 18464 9640 18528
rect 9704 18464 9710 18528
rect 9394 18463 9710 18464
rect 17842 18528 18158 18529
rect 17842 18464 17848 18528
rect 17912 18464 17928 18528
rect 17992 18464 18008 18528
rect 18072 18464 18088 18528
rect 18152 18464 18158 18528
rect 17842 18463 18158 18464
rect 26290 18528 26606 18529
rect 26290 18464 26296 18528
rect 26360 18464 26376 18528
rect 26440 18464 26456 18528
rect 26520 18464 26536 18528
rect 26600 18464 26606 18528
rect 26290 18463 26606 18464
rect 3417 18458 3483 18461
rect 0 18456 3483 18458
rect 0 18400 3422 18456
rect 3478 18400 3483 18456
rect 0 18398 3483 18400
rect 0 18308 800 18398
rect 3417 18395 3483 18398
rect 35200 18308 36000 18548
rect 5170 17984 5486 17985
rect 5170 17920 5176 17984
rect 5240 17920 5256 17984
rect 5320 17920 5336 17984
rect 5400 17920 5416 17984
rect 5480 17920 5486 17984
rect 5170 17919 5486 17920
rect 13618 17984 13934 17985
rect 13618 17920 13624 17984
rect 13688 17920 13704 17984
rect 13768 17920 13784 17984
rect 13848 17920 13864 17984
rect 13928 17920 13934 17984
rect 13618 17919 13934 17920
rect 22066 17984 22382 17985
rect 22066 17920 22072 17984
rect 22136 17920 22152 17984
rect 22216 17920 22232 17984
rect 22296 17920 22312 17984
rect 22376 17920 22382 17984
rect 22066 17919 22382 17920
rect 30514 17984 30830 17985
rect 30514 17920 30520 17984
rect 30584 17920 30600 17984
rect 30664 17920 30680 17984
rect 30744 17920 30760 17984
rect 30824 17920 30830 17984
rect 30514 17919 30830 17920
rect 0 17628 800 17868
rect 33041 17778 33107 17781
rect 35200 17778 36000 17868
rect 33041 17776 36000 17778
rect 33041 17720 33046 17776
rect 33102 17720 36000 17776
rect 33041 17718 36000 17720
rect 33041 17715 33107 17718
rect 35200 17628 36000 17718
rect 9394 17440 9710 17441
rect 9394 17376 9400 17440
rect 9464 17376 9480 17440
rect 9544 17376 9560 17440
rect 9624 17376 9640 17440
rect 9704 17376 9710 17440
rect 9394 17375 9710 17376
rect 17842 17440 18158 17441
rect 17842 17376 17848 17440
rect 17912 17376 17928 17440
rect 17992 17376 18008 17440
rect 18072 17376 18088 17440
rect 18152 17376 18158 17440
rect 17842 17375 18158 17376
rect 26290 17440 26606 17441
rect 26290 17376 26296 17440
rect 26360 17376 26376 17440
rect 26440 17376 26456 17440
rect 26520 17376 26536 17440
rect 26600 17376 26606 17440
rect 26290 17375 26606 17376
rect 0 17098 800 17188
rect 3233 17098 3299 17101
rect 0 17096 3299 17098
rect 0 17040 3238 17096
rect 3294 17040 3299 17096
rect 0 17038 3299 17040
rect 0 16948 800 17038
rect 3233 17035 3299 17038
rect 32305 17098 32371 17101
rect 35200 17098 36000 17188
rect 32305 17096 36000 17098
rect 32305 17040 32310 17096
rect 32366 17040 36000 17096
rect 32305 17038 36000 17040
rect 32305 17035 32371 17038
rect 35200 16948 36000 17038
rect 5170 16896 5486 16897
rect 5170 16832 5176 16896
rect 5240 16832 5256 16896
rect 5320 16832 5336 16896
rect 5400 16832 5416 16896
rect 5480 16832 5486 16896
rect 5170 16831 5486 16832
rect 13618 16896 13934 16897
rect 13618 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13784 16896
rect 13848 16832 13864 16896
rect 13928 16832 13934 16896
rect 13618 16831 13934 16832
rect 22066 16896 22382 16897
rect 22066 16832 22072 16896
rect 22136 16832 22152 16896
rect 22216 16832 22232 16896
rect 22296 16832 22312 16896
rect 22376 16832 22382 16896
rect 22066 16831 22382 16832
rect 30514 16896 30830 16897
rect 30514 16832 30520 16896
rect 30584 16832 30600 16896
rect 30664 16832 30680 16896
rect 30744 16832 30760 16896
rect 30824 16832 30830 16896
rect 30514 16831 30830 16832
rect 0 16268 800 16508
rect 34145 16418 34211 16421
rect 35200 16418 36000 16508
rect 34145 16416 36000 16418
rect 34145 16360 34150 16416
rect 34206 16360 36000 16416
rect 34145 16358 36000 16360
rect 34145 16355 34211 16358
rect 9394 16352 9710 16353
rect 9394 16288 9400 16352
rect 9464 16288 9480 16352
rect 9544 16288 9560 16352
rect 9624 16288 9640 16352
rect 9704 16288 9710 16352
rect 9394 16287 9710 16288
rect 17842 16352 18158 16353
rect 17842 16288 17848 16352
rect 17912 16288 17928 16352
rect 17992 16288 18008 16352
rect 18072 16288 18088 16352
rect 18152 16288 18158 16352
rect 17842 16287 18158 16288
rect 26290 16352 26606 16353
rect 26290 16288 26296 16352
rect 26360 16288 26376 16352
rect 26440 16288 26456 16352
rect 26520 16288 26536 16352
rect 26600 16288 26606 16352
rect 26290 16287 26606 16288
rect 35200 16268 36000 16358
rect 0 15738 800 15828
rect 5170 15808 5486 15809
rect 5170 15744 5176 15808
rect 5240 15744 5256 15808
rect 5320 15744 5336 15808
rect 5400 15744 5416 15808
rect 5480 15744 5486 15808
rect 5170 15743 5486 15744
rect 13618 15808 13934 15809
rect 13618 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13784 15808
rect 13848 15744 13864 15808
rect 13928 15744 13934 15808
rect 13618 15743 13934 15744
rect 22066 15808 22382 15809
rect 22066 15744 22072 15808
rect 22136 15744 22152 15808
rect 22216 15744 22232 15808
rect 22296 15744 22312 15808
rect 22376 15744 22382 15808
rect 22066 15743 22382 15744
rect 30514 15808 30830 15809
rect 30514 15744 30520 15808
rect 30584 15744 30600 15808
rect 30664 15744 30680 15808
rect 30744 15744 30760 15808
rect 30824 15744 30830 15808
rect 30514 15743 30830 15744
rect 4061 15738 4127 15741
rect 0 15736 4127 15738
rect 0 15680 4066 15736
rect 4122 15680 4127 15736
rect 0 15678 4127 15680
rect 0 15588 800 15678
rect 4061 15675 4127 15678
rect 35200 15588 36000 15828
rect 9394 15264 9710 15265
rect 9394 15200 9400 15264
rect 9464 15200 9480 15264
rect 9544 15200 9560 15264
rect 9624 15200 9640 15264
rect 9704 15200 9710 15264
rect 9394 15199 9710 15200
rect 17842 15264 18158 15265
rect 17842 15200 17848 15264
rect 17912 15200 17928 15264
rect 17992 15200 18008 15264
rect 18072 15200 18088 15264
rect 18152 15200 18158 15264
rect 17842 15199 18158 15200
rect 26290 15264 26606 15265
rect 26290 15200 26296 15264
rect 26360 15200 26376 15264
rect 26440 15200 26456 15264
rect 26520 15200 26536 15264
rect 26600 15200 26606 15264
rect 26290 15199 26606 15200
rect 0 14908 800 15148
rect 5170 14720 5486 14721
rect 5170 14656 5176 14720
rect 5240 14656 5256 14720
rect 5320 14656 5336 14720
rect 5400 14656 5416 14720
rect 5480 14656 5486 14720
rect 5170 14655 5486 14656
rect 13618 14720 13934 14721
rect 13618 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13784 14720
rect 13848 14656 13864 14720
rect 13928 14656 13934 14720
rect 13618 14655 13934 14656
rect 22066 14720 22382 14721
rect 22066 14656 22072 14720
rect 22136 14656 22152 14720
rect 22216 14656 22232 14720
rect 22296 14656 22312 14720
rect 22376 14656 22382 14720
rect 22066 14655 22382 14656
rect 30514 14720 30830 14721
rect 30514 14656 30520 14720
rect 30584 14656 30600 14720
rect 30664 14656 30680 14720
rect 30744 14656 30760 14720
rect 30824 14656 30830 14720
rect 30514 14655 30830 14656
rect 0 14378 800 14468
rect 1853 14378 1919 14381
rect 0 14376 1919 14378
rect 0 14320 1858 14376
rect 1914 14320 1919 14376
rect 0 14318 1919 14320
rect 0 14228 800 14318
rect 1853 14315 1919 14318
rect 31753 14378 31819 14381
rect 35200 14378 36000 14468
rect 31753 14376 36000 14378
rect 31753 14320 31758 14376
rect 31814 14320 36000 14376
rect 31753 14318 36000 14320
rect 31753 14315 31819 14318
rect 35200 14228 36000 14318
rect 9394 14176 9710 14177
rect 9394 14112 9400 14176
rect 9464 14112 9480 14176
rect 9544 14112 9560 14176
rect 9624 14112 9640 14176
rect 9704 14112 9710 14176
rect 9394 14111 9710 14112
rect 17842 14176 18158 14177
rect 17842 14112 17848 14176
rect 17912 14112 17928 14176
rect 17992 14112 18008 14176
rect 18072 14112 18088 14176
rect 18152 14112 18158 14176
rect 17842 14111 18158 14112
rect 26290 14176 26606 14177
rect 26290 14112 26296 14176
rect 26360 14112 26376 14176
rect 26440 14112 26456 14176
rect 26520 14112 26536 14176
rect 26600 14112 26606 14176
rect 26290 14111 26606 14112
rect 0 13698 800 13788
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13548 800 13638
rect 2773 13635 2839 13638
rect 32765 13698 32831 13701
rect 35200 13698 36000 13788
rect 32765 13696 36000 13698
rect 32765 13640 32770 13696
rect 32826 13640 36000 13696
rect 32765 13638 36000 13640
rect 32765 13635 32831 13638
rect 5170 13632 5486 13633
rect 5170 13568 5176 13632
rect 5240 13568 5256 13632
rect 5320 13568 5336 13632
rect 5400 13568 5416 13632
rect 5480 13568 5486 13632
rect 5170 13567 5486 13568
rect 13618 13632 13934 13633
rect 13618 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13784 13632
rect 13848 13568 13864 13632
rect 13928 13568 13934 13632
rect 13618 13567 13934 13568
rect 22066 13632 22382 13633
rect 22066 13568 22072 13632
rect 22136 13568 22152 13632
rect 22216 13568 22232 13632
rect 22296 13568 22312 13632
rect 22376 13568 22382 13632
rect 22066 13567 22382 13568
rect 30514 13632 30830 13633
rect 30514 13568 30520 13632
rect 30584 13568 30600 13632
rect 30664 13568 30680 13632
rect 30744 13568 30760 13632
rect 30824 13568 30830 13632
rect 30514 13567 30830 13568
rect 35200 13548 36000 13638
rect 9394 13088 9710 13089
rect 9394 13024 9400 13088
rect 9464 13024 9480 13088
rect 9544 13024 9560 13088
rect 9624 13024 9640 13088
rect 9704 13024 9710 13088
rect 9394 13023 9710 13024
rect 17842 13088 18158 13089
rect 17842 13024 17848 13088
rect 17912 13024 17928 13088
rect 17992 13024 18008 13088
rect 18072 13024 18088 13088
rect 18152 13024 18158 13088
rect 17842 13023 18158 13024
rect 26290 13088 26606 13089
rect 26290 13024 26296 13088
rect 26360 13024 26376 13088
rect 26440 13024 26456 13088
rect 26520 13024 26536 13088
rect 26600 13024 26606 13088
rect 26290 13023 26606 13024
rect 34145 13018 34211 13021
rect 35200 13018 36000 13108
rect 34145 13016 36000 13018
rect 34145 12960 34150 13016
rect 34206 12960 36000 13016
rect 34145 12958 36000 12960
rect 34145 12955 34211 12958
rect 35200 12868 36000 12958
rect 5170 12544 5486 12545
rect 5170 12480 5176 12544
rect 5240 12480 5256 12544
rect 5320 12480 5336 12544
rect 5400 12480 5416 12544
rect 5480 12480 5486 12544
rect 5170 12479 5486 12480
rect 13618 12544 13934 12545
rect 13618 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13784 12544
rect 13848 12480 13864 12544
rect 13928 12480 13934 12544
rect 13618 12479 13934 12480
rect 22066 12544 22382 12545
rect 22066 12480 22072 12544
rect 22136 12480 22152 12544
rect 22216 12480 22232 12544
rect 22296 12480 22312 12544
rect 22376 12480 22382 12544
rect 22066 12479 22382 12480
rect 30514 12544 30830 12545
rect 30514 12480 30520 12544
rect 30584 12480 30600 12544
rect 30664 12480 30680 12544
rect 30744 12480 30760 12544
rect 30824 12480 30830 12544
rect 30514 12479 30830 12480
rect 0 12188 800 12428
rect 33041 12338 33107 12341
rect 35200 12338 36000 12428
rect 33041 12336 36000 12338
rect 33041 12280 33046 12336
rect 33102 12280 36000 12336
rect 33041 12278 36000 12280
rect 33041 12275 33107 12278
rect 35200 12188 36000 12278
rect 9394 12000 9710 12001
rect 9394 11936 9400 12000
rect 9464 11936 9480 12000
rect 9544 11936 9560 12000
rect 9624 11936 9640 12000
rect 9704 11936 9710 12000
rect 9394 11935 9710 11936
rect 17842 12000 18158 12001
rect 17842 11936 17848 12000
rect 17912 11936 17928 12000
rect 17992 11936 18008 12000
rect 18072 11936 18088 12000
rect 18152 11936 18158 12000
rect 17842 11935 18158 11936
rect 26290 12000 26606 12001
rect 26290 11936 26296 12000
rect 26360 11936 26376 12000
rect 26440 11936 26456 12000
rect 26520 11936 26536 12000
rect 26600 11936 26606 12000
rect 26290 11935 26606 11936
rect 0 11658 800 11748
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11508 800 11598
rect 4061 11595 4127 11598
rect 35200 11508 36000 11748
rect 5170 11456 5486 11457
rect 5170 11392 5176 11456
rect 5240 11392 5256 11456
rect 5320 11392 5336 11456
rect 5400 11392 5416 11456
rect 5480 11392 5486 11456
rect 5170 11391 5486 11392
rect 13618 11456 13934 11457
rect 13618 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13784 11456
rect 13848 11392 13864 11456
rect 13928 11392 13934 11456
rect 13618 11391 13934 11392
rect 22066 11456 22382 11457
rect 22066 11392 22072 11456
rect 22136 11392 22152 11456
rect 22216 11392 22232 11456
rect 22296 11392 22312 11456
rect 22376 11392 22382 11456
rect 22066 11391 22382 11392
rect 30514 11456 30830 11457
rect 30514 11392 30520 11456
rect 30584 11392 30600 11456
rect 30664 11392 30680 11456
rect 30744 11392 30760 11456
rect 30824 11392 30830 11456
rect 30514 11391 30830 11392
rect 0 10978 800 11068
rect 2773 10978 2839 10981
rect 0 10976 2839 10978
rect 0 10920 2778 10976
rect 2834 10920 2839 10976
rect 0 10918 2839 10920
rect 0 10828 800 10918
rect 2773 10915 2839 10918
rect 9394 10912 9710 10913
rect 9394 10848 9400 10912
rect 9464 10848 9480 10912
rect 9544 10848 9560 10912
rect 9624 10848 9640 10912
rect 9704 10848 9710 10912
rect 9394 10847 9710 10848
rect 17842 10912 18158 10913
rect 17842 10848 17848 10912
rect 17912 10848 17928 10912
rect 17992 10848 18008 10912
rect 18072 10848 18088 10912
rect 18152 10848 18158 10912
rect 17842 10847 18158 10848
rect 26290 10912 26606 10913
rect 26290 10848 26296 10912
rect 26360 10848 26376 10912
rect 26440 10848 26456 10912
rect 26520 10848 26536 10912
rect 26600 10848 26606 10912
rect 26290 10847 26606 10848
rect 35200 10828 36000 11068
rect 0 10148 800 10388
rect 5170 10368 5486 10369
rect 5170 10304 5176 10368
rect 5240 10304 5256 10368
rect 5320 10304 5336 10368
rect 5400 10304 5416 10368
rect 5480 10304 5486 10368
rect 5170 10303 5486 10304
rect 13618 10368 13934 10369
rect 13618 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13784 10368
rect 13848 10304 13864 10368
rect 13928 10304 13934 10368
rect 13618 10303 13934 10304
rect 22066 10368 22382 10369
rect 22066 10304 22072 10368
rect 22136 10304 22152 10368
rect 22216 10304 22232 10368
rect 22296 10304 22312 10368
rect 22376 10304 22382 10368
rect 22066 10303 22382 10304
rect 30514 10368 30830 10369
rect 30514 10304 30520 10368
rect 30584 10304 30600 10368
rect 30664 10304 30680 10368
rect 30744 10304 30760 10368
rect 30824 10304 30830 10368
rect 30514 10303 30830 10304
rect 35200 10148 36000 10388
rect 9394 9824 9710 9825
rect 9394 9760 9400 9824
rect 9464 9760 9480 9824
rect 9544 9760 9560 9824
rect 9624 9760 9640 9824
rect 9704 9760 9710 9824
rect 9394 9759 9710 9760
rect 17842 9824 18158 9825
rect 17842 9760 17848 9824
rect 17912 9760 17928 9824
rect 17992 9760 18008 9824
rect 18072 9760 18088 9824
rect 18152 9760 18158 9824
rect 17842 9759 18158 9760
rect 26290 9824 26606 9825
rect 26290 9760 26296 9824
rect 26360 9760 26376 9824
rect 26440 9760 26456 9824
rect 26520 9760 26536 9824
rect 26600 9760 26606 9824
rect 26290 9759 26606 9760
rect 0 9468 800 9708
rect 35200 9468 36000 9708
rect 5170 9280 5486 9281
rect 5170 9216 5176 9280
rect 5240 9216 5256 9280
rect 5320 9216 5336 9280
rect 5400 9216 5416 9280
rect 5480 9216 5486 9280
rect 5170 9215 5486 9216
rect 13618 9280 13934 9281
rect 13618 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13784 9280
rect 13848 9216 13864 9280
rect 13928 9216 13934 9280
rect 13618 9215 13934 9216
rect 22066 9280 22382 9281
rect 22066 9216 22072 9280
rect 22136 9216 22152 9280
rect 22216 9216 22232 9280
rect 22296 9216 22312 9280
rect 22376 9216 22382 9280
rect 22066 9215 22382 9216
rect 30514 9280 30830 9281
rect 30514 9216 30520 9280
rect 30584 9216 30600 9280
rect 30664 9216 30680 9280
rect 30744 9216 30760 9280
rect 30824 9216 30830 9280
rect 30514 9215 30830 9216
rect 0 8938 800 9028
rect 1853 8938 1919 8941
rect 0 8936 1919 8938
rect 0 8880 1858 8936
rect 1914 8880 1919 8936
rect 0 8878 1919 8880
rect 0 8788 800 8878
rect 1853 8875 1919 8878
rect 31753 8938 31819 8941
rect 35200 8938 36000 9028
rect 31753 8936 36000 8938
rect 31753 8880 31758 8936
rect 31814 8880 36000 8936
rect 31753 8878 36000 8880
rect 31753 8875 31819 8878
rect 35200 8788 36000 8878
rect 9394 8736 9710 8737
rect 9394 8672 9400 8736
rect 9464 8672 9480 8736
rect 9544 8672 9560 8736
rect 9624 8672 9640 8736
rect 9704 8672 9710 8736
rect 9394 8671 9710 8672
rect 17842 8736 18158 8737
rect 17842 8672 17848 8736
rect 17912 8672 17928 8736
rect 17992 8672 18008 8736
rect 18072 8672 18088 8736
rect 18152 8672 18158 8736
rect 17842 8671 18158 8672
rect 26290 8736 26606 8737
rect 26290 8672 26296 8736
rect 26360 8672 26376 8736
rect 26440 8672 26456 8736
rect 26520 8672 26536 8736
rect 26600 8672 26606 8736
rect 26290 8671 26606 8672
rect 0 8258 800 8348
rect 3141 8258 3207 8261
rect 0 8256 3207 8258
rect 0 8200 3146 8256
rect 3202 8200 3207 8256
rect 0 8198 3207 8200
rect 0 8108 800 8198
rect 3141 8195 3207 8198
rect 5170 8192 5486 8193
rect 5170 8128 5176 8192
rect 5240 8128 5256 8192
rect 5320 8128 5336 8192
rect 5400 8128 5416 8192
rect 5480 8128 5486 8192
rect 5170 8127 5486 8128
rect 13618 8192 13934 8193
rect 13618 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13784 8192
rect 13848 8128 13864 8192
rect 13928 8128 13934 8192
rect 13618 8127 13934 8128
rect 22066 8192 22382 8193
rect 22066 8128 22072 8192
rect 22136 8128 22152 8192
rect 22216 8128 22232 8192
rect 22296 8128 22312 8192
rect 22376 8128 22382 8192
rect 22066 8127 22382 8128
rect 30514 8192 30830 8193
rect 30514 8128 30520 8192
rect 30584 8128 30600 8192
rect 30664 8128 30680 8192
rect 30744 8128 30760 8192
rect 30824 8128 30830 8192
rect 30514 8127 30830 8128
rect 0 7578 800 7668
rect 9394 7648 9710 7649
rect 9394 7584 9400 7648
rect 9464 7584 9480 7648
rect 9544 7584 9560 7648
rect 9624 7584 9640 7648
rect 9704 7584 9710 7648
rect 9394 7583 9710 7584
rect 17842 7648 18158 7649
rect 17842 7584 17848 7648
rect 17912 7584 17928 7648
rect 17992 7584 18008 7648
rect 18072 7584 18088 7648
rect 18152 7584 18158 7648
rect 17842 7583 18158 7584
rect 26290 7648 26606 7649
rect 26290 7584 26296 7648
rect 26360 7584 26376 7648
rect 26440 7584 26456 7648
rect 26520 7584 26536 7648
rect 26600 7584 26606 7648
rect 26290 7583 26606 7584
rect 3141 7578 3207 7581
rect 0 7576 3207 7578
rect 0 7520 3146 7576
rect 3202 7520 3207 7576
rect 0 7518 3207 7520
rect 0 7428 800 7518
rect 3141 7515 3207 7518
rect 35200 7428 36000 7668
rect 5170 7104 5486 7105
rect 5170 7040 5176 7104
rect 5240 7040 5256 7104
rect 5320 7040 5336 7104
rect 5400 7040 5416 7104
rect 5480 7040 5486 7104
rect 5170 7039 5486 7040
rect 13618 7104 13934 7105
rect 13618 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13784 7104
rect 13848 7040 13864 7104
rect 13928 7040 13934 7104
rect 13618 7039 13934 7040
rect 22066 7104 22382 7105
rect 22066 7040 22072 7104
rect 22136 7040 22152 7104
rect 22216 7040 22232 7104
rect 22296 7040 22312 7104
rect 22376 7040 22382 7104
rect 22066 7039 22382 7040
rect 30514 7104 30830 7105
rect 30514 7040 30520 7104
rect 30584 7040 30600 7104
rect 30664 7040 30680 7104
rect 30744 7040 30760 7104
rect 30824 7040 30830 7104
rect 30514 7039 30830 7040
rect 0 6748 800 6988
rect 34145 6898 34211 6901
rect 35200 6898 36000 6988
rect 34145 6896 36000 6898
rect 34145 6840 34150 6896
rect 34206 6840 36000 6896
rect 34145 6838 36000 6840
rect 34145 6835 34211 6838
rect 35200 6748 36000 6838
rect 9394 6560 9710 6561
rect 9394 6496 9400 6560
rect 9464 6496 9480 6560
rect 9544 6496 9560 6560
rect 9624 6496 9640 6560
rect 9704 6496 9710 6560
rect 9394 6495 9710 6496
rect 17842 6560 18158 6561
rect 17842 6496 17848 6560
rect 17912 6496 17928 6560
rect 17992 6496 18008 6560
rect 18072 6496 18088 6560
rect 18152 6496 18158 6560
rect 17842 6495 18158 6496
rect 26290 6560 26606 6561
rect 26290 6496 26296 6560
rect 26360 6496 26376 6560
rect 26440 6496 26456 6560
rect 26520 6496 26536 6560
rect 26600 6496 26606 6560
rect 26290 6495 26606 6496
rect 35200 6068 36000 6308
rect 5170 6016 5486 6017
rect 5170 5952 5176 6016
rect 5240 5952 5256 6016
rect 5320 5952 5336 6016
rect 5400 5952 5416 6016
rect 5480 5952 5486 6016
rect 5170 5951 5486 5952
rect 13618 6016 13934 6017
rect 13618 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13784 6016
rect 13848 5952 13864 6016
rect 13928 5952 13934 6016
rect 13618 5951 13934 5952
rect 22066 6016 22382 6017
rect 22066 5952 22072 6016
rect 22136 5952 22152 6016
rect 22216 5952 22232 6016
rect 22296 5952 22312 6016
rect 22376 5952 22382 6016
rect 22066 5951 22382 5952
rect 30514 6016 30830 6017
rect 30514 5952 30520 6016
rect 30584 5952 30600 6016
rect 30664 5952 30680 6016
rect 30744 5952 30760 6016
rect 30824 5952 30830 6016
rect 30514 5951 30830 5952
rect 0 5538 800 5628
rect 3417 5538 3483 5541
rect 0 5536 3483 5538
rect 0 5480 3422 5536
rect 3478 5480 3483 5536
rect 0 5478 3483 5480
rect 0 5388 800 5478
rect 3417 5475 3483 5478
rect 9394 5472 9710 5473
rect 9394 5408 9400 5472
rect 9464 5408 9480 5472
rect 9544 5408 9560 5472
rect 9624 5408 9640 5472
rect 9704 5408 9710 5472
rect 9394 5407 9710 5408
rect 17842 5472 18158 5473
rect 17842 5408 17848 5472
rect 17912 5408 17928 5472
rect 17992 5408 18008 5472
rect 18072 5408 18088 5472
rect 18152 5408 18158 5472
rect 17842 5407 18158 5408
rect 26290 5472 26606 5473
rect 26290 5408 26296 5472
rect 26360 5408 26376 5472
rect 26440 5408 26456 5472
rect 26520 5408 26536 5472
rect 26600 5408 26606 5472
rect 26290 5407 26606 5408
rect 35200 5388 36000 5628
rect 0 4858 800 4948
rect 5170 4928 5486 4929
rect 5170 4864 5176 4928
rect 5240 4864 5256 4928
rect 5320 4864 5336 4928
rect 5400 4864 5416 4928
rect 5480 4864 5486 4928
rect 5170 4863 5486 4864
rect 13618 4928 13934 4929
rect 13618 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13784 4928
rect 13848 4864 13864 4928
rect 13928 4864 13934 4928
rect 13618 4863 13934 4864
rect 22066 4928 22382 4929
rect 22066 4864 22072 4928
rect 22136 4864 22152 4928
rect 22216 4864 22232 4928
rect 22296 4864 22312 4928
rect 22376 4864 22382 4928
rect 22066 4863 22382 4864
rect 30514 4928 30830 4929
rect 30514 4864 30520 4928
rect 30584 4864 30600 4928
rect 30664 4864 30680 4928
rect 30744 4864 30760 4928
rect 30824 4864 30830 4928
rect 30514 4863 30830 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4708 800 4798
rect 2773 4795 2839 4798
rect 32305 4858 32371 4861
rect 35200 4858 36000 4948
rect 32305 4856 36000 4858
rect 32305 4800 32310 4856
rect 32366 4800 36000 4856
rect 32305 4798 36000 4800
rect 32305 4795 32371 4798
rect 35200 4708 36000 4798
rect 9394 4384 9710 4385
rect 9394 4320 9400 4384
rect 9464 4320 9480 4384
rect 9544 4320 9560 4384
rect 9624 4320 9640 4384
rect 9704 4320 9710 4384
rect 9394 4319 9710 4320
rect 17842 4384 18158 4385
rect 17842 4320 17848 4384
rect 17912 4320 17928 4384
rect 17992 4320 18008 4384
rect 18072 4320 18088 4384
rect 18152 4320 18158 4384
rect 17842 4319 18158 4320
rect 26290 4384 26606 4385
rect 26290 4320 26296 4384
rect 26360 4320 26376 4384
rect 26440 4320 26456 4384
rect 26520 4320 26536 4384
rect 26600 4320 26606 4384
rect 26290 4319 26606 4320
rect 0 4178 800 4268
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4028 800 4118
rect 3417 4115 3483 4118
rect 32397 4178 32463 4181
rect 35200 4178 36000 4268
rect 32397 4176 36000 4178
rect 32397 4120 32402 4176
rect 32458 4120 36000 4176
rect 32397 4118 36000 4120
rect 32397 4115 32463 4118
rect 35200 4028 36000 4118
rect 5170 3840 5486 3841
rect 5170 3776 5176 3840
rect 5240 3776 5256 3840
rect 5320 3776 5336 3840
rect 5400 3776 5416 3840
rect 5480 3776 5486 3840
rect 5170 3775 5486 3776
rect 13618 3840 13934 3841
rect 13618 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13784 3840
rect 13848 3776 13864 3840
rect 13928 3776 13934 3840
rect 13618 3775 13934 3776
rect 22066 3840 22382 3841
rect 22066 3776 22072 3840
rect 22136 3776 22152 3840
rect 22216 3776 22232 3840
rect 22296 3776 22312 3840
rect 22376 3776 22382 3840
rect 22066 3775 22382 3776
rect 30514 3840 30830 3841
rect 30514 3776 30520 3840
rect 30584 3776 30600 3840
rect 30664 3776 30680 3840
rect 30744 3776 30760 3840
rect 30824 3776 30830 3840
rect 30514 3775 30830 3776
rect 0 3498 800 3588
rect 3417 3498 3483 3501
rect 0 3496 3483 3498
rect 0 3440 3422 3496
rect 3478 3440 3483 3496
rect 0 3438 3483 3440
rect 0 3348 800 3438
rect 3417 3435 3483 3438
rect 33041 3498 33107 3501
rect 35200 3498 36000 3588
rect 33041 3496 36000 3498
rect 33041 3440 33046 3496
rect 33102 3440 36000 3496
rect 33041 3438 36000 3440
rect 33041 3435 33107 3438
rect 35200 3348 36000 3438
rect 9394 3296 9710 3297
rect 9394 3232 9400 3296
rect 9464 3232 9480 3296
rect 9544 3232 9560 3296
rect 9624 3232 9640 3296
rect 9704 3232 9710 3296
rect 9394 3231 9710 3232
rect 17842 3296 18158 3297
rect 17842 3232 17848 3296
rect 17912 3232 17928 3296
rect 17992 3232 18008 3296
rect 18072 3232 18088 3296
rect 18152 3232 18158 3296
rect 17842 3231 18158 3232
rect 26290 3296 26606 3297
rect 26290 3232 26296 3296
rect 26360 3232 26376 3296
rect 26440 3232 26456 3296
rect 26520 3232 26536 3296
rect 26600 3232 26606 3296
rect 26290 3231 26606 3232
rect 0 2818 800 2908
rect 3417 2818 3483 2821
rect 0 2816 3483 2818
rect 0 2760 3422 2816
rect 3478 2760 3483 2816
rect 0 2758 3483 2760
rect 0 2668 800 2758
rect 3417 2755 3483 2758
rect 5170 2752 5486 2753
rect 5170 2688 5176 2752
rect 5240 2688 5256 2752
rect 5320 2688 5336 2752
rect 5400 2688 5416 2752
rect 5480 2688 5486 2752
rect 5170 2687 5486 2688
rect 13618 2752 13934 2753
rect 13618 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13784 2752
rect 13848 2688 13864 2752
rect 13928 2688 13934 2752
rect 13618 2687 13934 2688
rect 22066 2752 22382 2753
rect 22066 2688 22072 2752
rect 22136 2688 22152 2752
rect 22216 2688 22232 2752
rect 22296 2688 22312 2752
rect 22376 2688 22382 2752
rect 22066 2687 22382 2688
rect 30514 2752 30830 2753
rect 30514 2688 30520 2752
rect 30584 2688 30600 2752
rect 30664 2688 30680 2752
rect 30744 2688 30760 2752
rect 30824 2688 30830 2752
rect 30514 2687 30830 2688
rect 35200 2668 36000 2908
rect 0 2138 800 2228
rect 9394 2208 9710 2209
rect 9394 2144 9400 2208
rect 9464 2144 9480 2208
rect 9544 2144 9560 2208
rect 9624 2144 9640 2208
rect 9704 2144 9710 2208
rect 9394 2143 9710 2144
rect 17842 2208 18158 2209
rect 17842 2144 17848 2208
rect 17912 2144 17928 2208
rect 17992 2144 18008 2208
rect 18072 2144 18088 2208
rect 18152 2144 18158 2208
rect 17842 2143 18158 2144
rect 26290 2208 26606 2209
rect 26290 2144 26296 2208
rect 26360 2144 26376 2208
rect 26440 2144 26456 2208
rect 26520 2144 26536 2208
rect 26600 2144 26606 2208
rect 26290 2143 26606 2144
rect 3417 2138 3483 2141
rect 0 2136 3483 2138
rect 0 2080 3422 2136
rect 3478 2080 3483 2136
rect 0 2078 3483 2080
rect 0 1988 800 2078
rect 3417 2075 3483 2078
rect 31753 2138 31819 2141
rect 35200 2138 36000 2228
rect 31753 2136 36000 2138
rect 31753 2080 31758 2136
rect 31814 2080 36000 2136
rect 31753 2078 36000 2080
rect 31753 2075 31819 2078
rect 35200 1988 36000 2078
rect 0 1458 800 1548
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1308 800 1398
rect 3325 1395 3391 1398
rect 0 628 800 868
rect 31385 778 31451 781
rect 35200 778 36000 868
rect 31385 776 36000 778
rect 31385 720 31390 776
rect 31446 720 36000 776
rect 31385 718 36000 720
rect 31385 715 31451 718
rect 35200 628 36000 718
rect 33961 98 34027 101
rect 35200 98 36000 188
rect 33961 96 36000 98
rect 33961 40 33966 96
rect 34022 40 36000 96
rect 33961 38 36000 40
rect 33961 35 34027 38
rect 35200 -52 36000 38
<< via3 >>
rect 5176 39740 5240 39744
rect 5176 39684 5180 39740
rect 5180 39684 5236 39740
rect 5236 39684 5240 39740
rect 5176 39680 5240 39684
rect 5256 39740 5320 39744
rect 5256 39684 5260 39740
rect 5260 39684 5316 39740
rect 5316 39684 5320 39740
rect 5256 39680 5320 39684
rect 5336 39740 5400 39744
rect 5336 39684 5340 39740
rect 5340 39684 5396 39740
rect 5396 39684 5400 39740
rect 5336 39680 5400 39684
rect 5416 39740 5480 39744
rect 5416 39684 5420 39740
rect 5420 39684 5476 39740
rect 5476 39684 5480 39740
rect 5416 39680 5480 39684
rect 13624 39740 13688 39744
rect 13624 39684 13628 39740
rect 13628 39684 13684 39740
rect 13684 39684 13688 39740
rect 13624 39680 13688 39684
rect 13704 39740 13768 39744
rect 13704 39684 13708 39740
rect 13708 39684 13764 39740
rect 13764 39684 13768 39740
rect 13704 39680 13768 39684
rect 13784 39740 13848 39744
rect 13784 39684 13788 39740
rect 13788 39684 13844 39740
rect 13844 39684 13848 39740
rect 13784 39680 13848 39684
rect 13864 39740 13928 39744
rect 13864 39684 13868 39740
rect 13868 39684 13924 39740
rect 13924 39684 13928 39740
rect 13864 39680 13928 39684
rect 22072 39740 22136 39744
rect 22072 39684 22076 39740
rect 22076 39684 22132 39740
rect 22132 39684 22136 39740
rect 22072 39680 22136 39684
rect 22152 39740 22216 39744
rect 22152 39684 22156 39740
rect 22156 39684 22212 39740
rect 22212 39684 22216 39740
rect 22152 39680 22216 39684
rect 22232 39740 22296 39744
rect 22232 39684 22236 39740
rect 22236 39684 22292 39740
rect 22292 39684 22296 39740
rect 22232 39680 22296 39684
rect 22312 39740 22376 39744
rect 22312 39684 22316 39740
rect 22316 39684 22372 39740
rect 22372 39684 22376 39740
rect 22312 39680 22376 39684
rect 30520 39740 30584 39744
rect 30520 39684 30524 39740
rect 30524 39684 30580 39740
rect 30580 39684 30584 39740
rect 30520 39680 30584 39684
rect 30600 39740 30664 39744
rect 30600 39684 30604 39740
rect 30604 39684 30660 39740
rect 30660 39684 30664 39740
rect 30600 39680 30664 39684
rect 30680 39740 30744 39744
rect 30680 39684 30684 39740
rect 30684 39684 30740 39740
rect 30740 39684 30744 39740
rect 30680 39680 30744 39684
rect 30760 39740 30824 39744
rect 30760 39684 30764 39740
rect 30764 39684 30820 39740
rect 30820 39684 30824 39740
rect 30760 39680 30824 39684
rect 9400 39196 9464 39200
rect 9400 39140 9404 39196
rect 9404 39140 9460 39196
rect 9460 39140 9464 39196
rect 9400 39136 9464 39140
rect 9480 39196 9544 39200
rect 9480 39140 9484 39196
rect 9484 39140 9540 39196
rect 9540 39140 9544 39196
rect 9480 39136 9544 39140
rect 9560 39196 9624 39200
rect 9560 39140 9564 39196
rect 9564 39140 9620 39196
rect 9620 39140 9624 39196
rect 9560 39136 9624 39140
rect 9640 39196 9704 39200
rect 9640 39140 9644 39196
rect 9644 39140 9700 39196
rect 9700 39140 9704 39196
rect 9640 39136 9704 39140
rect 17848 39196 17912 39200
rect 17848 39140 17852 39196
rect 17852 39140 17908 39196
rect 17908 39140 17912 39196
rect 17848 39136 17912 39140
rect 17928 39196 17992 39200
rect 17928 39140 17932 39196
rect 17932 39140 17988 39196
rect 17988 39140 17992 39196
rect 17928 39136 17992 39140
rect 18008 39196 18072 39200
rect 18008 39140 18012 39196
rect 18012 39140 18068 39196
rect 18068 39140 18072 39196
rect 18008 39136 18072 39140
rect 18088 39196 18152 39200
rect 18088 39140 18092 39196
rect 18092 39140 18148 39196
rect 18148 39140 18152 39196
rect 18088 39136 18152 39140
rect 26296 39196 26360 39200
rect 26296 39140 26300 39196
rect 26300 39140 26356 39196
rect 26356 39140 26360 39196
rect 26296 39136 26360 39140
rect 26376 39196 26440 39200
rect 26376 39140 26380 39196
rect 26380 39140 26436 39196
rect 26436 39140 26440 39196
rect 26376 39136 26440 39140
rect 26456 39196 26520 39200
rect 26456 39140 26460 39196
rect 26460 39140 26516 39196
rect 26516 39140 26520 39196
rect 26456 39136 26520 39140
rect 26536 39196 26600 39200
rect 26536 39140 26540 39196
rect 26540 39140 26596 39196
rect 26596 39140 26600 39196
rect 26536 39136 26600 39140
rect 5176 38652 5240 38656
rect 5176 38596 5180 38652
rect 5180 38596 5236 38652
rect 5236 38596 5240 38652
rect 5176 38592 5240 38596
rect 5256 38652 5320 38656
rect 5256 38596 5260 38652
rect 5260 38596 5316 38652
rect 5316 38596 5320 38652
rect 5256 38592 5320 38596
rect 5336 38652 5400 38656
rect 5336 38596 5340 38652
rect 5340 38596 5396 38652
rect 5396 38596 5400 38652
rect 5336 38592 5400 38596
rect 5416 38652 5480 38656
rect 5416 38596 5420 38652
rect 5420 38596 5476 38652
rect 5476 38596 5480 38652
rect 5416 38592 5480 38596
rect 13624 38652 13688 38656
rect 13624 38596 13628 38652
rect 13628 38596 13684 38652
rect 13684 38596 13688 38652
rect 13624 38592 13688 38596
rect 13704 38652 13768 38656
rect 13704 38596 13708 38652
rect 13708 38596 13764 38652
rect 13764 38596 13768 38652
rect 13704 38592 13768 38596
rect 13784 38652 13848 38656
rect 13784 38596 13788 38652
rect 13788 38596 13844 38652
rect 13844 38596 13848 38652
rect 13784 38592 13848 38596
rect 13864 38652 13928 38656
rect 13864 38596 13868 38652
rect 13868 38596 13924 38652
rect 13924 38596 13928 38652
rect 13864 38592 13928 38596
rect 22072 38652 22136 38656
rect 22072 38596 22076 38652
rect 22076 38596 22132 38652
rect 22132 38596 22136 38652
rect 22072 38592 22136 38596
rect 22152 38652 22216 38656
rect 22152 38596 22156 38652
rect 22156 38596 22212 38652
rect 22212 38596 22216 38652
rect 22152 38592 22216 38596
rect 22232 38652 22296 38656
rect 22232 38596 22236 38652
rect 22236 38596 22292 38652
rect 22292 38596 22296 38652
rect 22232 38592 22296 38596
rect 22312 38652 22376 38656
rect 22312 38596 22316 38652
rect 22316 38596 22372 38652
rect 22372 38596 22376 38652
rect 22312 38592 22376 38596
rect 30520 38652 30584 38656
rect 30520 38596 30524 38652
rect 30524 38596 30580 38652
rect 30580 38596 30584 38652
rect 30520 38592 30584 38596
rect 30600 38652 30664 38656
rect 30600 38596 30604 38652
rect 30604 38596 30660 38652
rect 30660 38596 30664 38652
rect 30600 38592 30664 38596
rect 30680 38652 30744 38656
rect 30680 38596 30684 38652
rect 30684 38596 30740 38652
rect 30740 38596 30744 38652
rect 30680 38592 30744 38596
rect 30760 38652 30824 38656
rect 30760 38596 30764 38652
rect 30764 38596 30820 38652
rect 30820 38596 30824 38652
rect 30760 38592 30824 38596
rect 9400 38108 9464 38112
rect 9400 38052 9404 38108
rect 9404 38052 9460 38108
rect 9460 38052 9464 38108
rect 9400 38048 9464 38052
rect 9480 38108 9544 38112
rect 9480 38052 9484 38108
rect 9484 38052 9540 38108
rect 9540 38052 9544 38108
rect 9480 38048 9544 38052
rect 9560 38108 9624 38112
rect 9560 38052 9564 38108
rect 9564 38052 9620 38108
rect 9620 38052 9624 38108
rect 9560 38048 9624 38052
rect 9640 38108 9704 38112
rect 9640 38052 9644 38108
rect 9644 38052 9700 38108
rect 9700 38052 9704 38108
rect 9640 38048 9704 38052
rect 17848 38108 17912 38112
rect 17848 38052 17852 38108
rect 17852 38052 17908 38108
rect 17908 38052 17912 38108
rect 17848 38048 17912 38052
rect 17928 38108 17992 38112
rect 17928 38052 17932 38108
rect 17932 38052 17988 38108
rect 17988 38052 17992 38108
rect 17928 38048 17992 38052
rect 18008 38108 18072 38112
rect 18008 38052 18012 38108
rect 18012 38052 18068 38108
rect 18068 38052 18072 38108
rect 18008 38048 18072 38052
rect 18088 38108 18152 38112
rect 18088 38052 18092 38108
rect 18092 38052 18148 38108
rect 18148 38052 18152 38108
rect 18088 38048 18152 38052
rect 26296 38108 26360 38112
rect 26296 38052 26300 38108
rect 26300 38052 26356 38108
rect 26356 38052 26360 38108
rect 26296 38048 26360 38052
rect 26376 38108 26440 38112
rect 26376 38052 26380 38108
rect 26380 38052 26436 38108
rect 26436 38052 26440 38108
rect 26376 38048 26440 38052
rect 26456 38108 26520 38112
rect 26456 38052 26460 38108
rect 26460 38052 26516 38108
rect 26516 38052 26520 38108
rect 26456 38048 26520 38052
rect 26536 38108 26600 38112
rect 26536 38052 26540 38108
rect 26540 38052 26596 38108
rect 26596 38052 26600 38108
rect 26536 38048 26600 38052
rect 5176 37564 5240 37568
rect 5176 37508 5180 37564
rect 5180 37508 5236 37564
rect 5236 37508 5240 37564
rect 5176 37504 5240 37508
rect 5256 37564 5320 37568
rect 5256 37508 5260 37564
rect 5260 37508 5316 37564
rect 5316 37508 5320 37564
rect 5256 37504 5320 37508
rect 5336 37564 5400 37568
rect 5336 37508 5340 37564
rect 5340 37508 5396 37564
rect 5396 37508 5400 37564
rect 5336 37504 5400 37508
rect 5416 37564 5480 37568
rect 5416 37508 5420 37564
rect 5420 37508 5476 37564
rect 5476 37508 5480 37564
rect 5416 37504 5480 37508
rect 13624 37564 13688 37568
rect 13624 37508 13628 37564
rect 13628 37508 13684 37564
rect 13684 37508 13688 37564
rect 13624 37504 13688 37508
rect 13704 37564 13768 37568
rect 13704 37508 13708 37564
rect 13708 37508 13764 37564
rect 13764 37508 13768 37564
rect 13704 37504 13768 37508
rect 13784 37564 13848 37568
rect 13784 37508 13788 37564
rect 13788 37508 13844 37564
rect 13844 37508 13848 37564
rect 13784 37504 13848 37508
rect 13864 37564 13928 37568
rect 13864 37508 13868 37564
rect 13868 37508 13924 37564
rect 13924 37508 13928 37564
rect 13864 37504 13928 37508
rect 22072 37564 22136 37568
rect 22072 37508 22076 37564
rect 22076 37508 22132 37564
rect 22132 37508 22136 37564
rect 22072 37504 22136 37508
rect 22152 37564 22216 37568
rect 22152 37508 22156 37564
rect 22156 37508 22212 37564
rect 22212 37508 22216 37564
rect 22152 37504 22216 37508
rect 22232 37564 22296 37568
rect 22232 37508 22236 37564
rect 22236 37508 22292 37564
rect 22292 37508 22296 37564
rect 22232 37504 22296 37508
rect 22312 37564 22376 37568
rect 22312 37508 22316 37564
rect 22316 37508 22372 37564
rect 22372 37508 22376 37564
rect 22312 37504 22376 37508
rect 30520 37564 30584 37568
rect 30520 37508 30524 37564
rect 30524 37508 30580 37564
rect 30580 37508 30584 37564
rect 30520 37504 30584 37508
rect 30600 37564 30664 37568
rect 30600 37508 30604 37564
rect 30604 37508 30660 37564
rect 30660 37508 30664 37564
rect 30600 37504 30664 37508
rect 30680 37564 30744 37568
rect 30680 37508 30684 37564
rect 30684 37508 30740 37564
rect 30740 37508 30744 37564
rect 30680 37504 30744 37508
rect 30760 37564 30824 37568
rect 30760 37508 30764 37564
rect 30764 37508 30820 37564
rect 30820 37508 30824 37564
rect 30760 37504 30824 37508
rect 9400 37020 9464 37024
rect 9400 36964 9404 37020
rect 9404 36964 9460 37020
rect 9460 36964 9464 37020
rect 9400 36960 9464 36964
rect 9480 37020 9544 37024
rect 9480 36964 9484 37020
rect 9484 36964 9540 37020
rect 9540 36964 9544 37020
rect 9480 36960 9544 36964
rect 9560 37020 9624 37024
rect 9560 36964 9564 37020
rect 9564 36964 9620 37020
rect 9620 36964 9624 37020
rect 9560 36960 9624 36964
rect 9640 37020 9704 37024
rect 9640 36964 9644 37020
rect 9644 36964 9700 37020
rect 9700 36964 9704 37020
rect 9640 36960 9704 36964
rect 17848 37020 17912 37024
rect 17848 36964 17852 37020
rect 17852 36964 17908 37020
rect 17908 36964 17912 37020
rect 17848 36960 17912 36964
rect 17928 37020 17992 37024
rect 17928 36964 17932 37020
rect 17932 36964 17988 37020
rect 17988 36964 17992 37020
rect 17928 36960 17992 36964
rect 18008 37020 18072 37024
rect 18008 36964 18012 37020
rect 18012 36964 18068 37020
rect 18068 36964 18072 37020
rect 18008 36960 18072 36964
rect 18088 37020 18152 37024
rect 18088 36964 18092 37020
rect 18092 36964 18148 37020
rect 18148 36964 18152 37020
rect 18088 36960 18152 36964
rect 26296 37020 26360 37024
rect 26296 36964 26300 37020
rect 26300 36964 26356 37020
rect 26356 36964 26360 37020
rect 26296 36960 26360 36964
rect 26376 37020 26440 37024
rect 26376 36964 26380 37020
rect 26380 36964 26436 37020
rect 26436 36964 26440 37020
rect 26376 36960 26440 36964
rect 26456 37020 26520 37024
rect 26456 36964 26460 37020
rect 26460 36964 26516 37020
rect 26516 36964 26520 37020
rect 26456 36960 26520 36964
rect 26536 37020 26600 37024
rect 26536 36964 26540 37020
rect 26540 36964 26596 37020
rect 26596 36964 26600 37020
rect 26536 36960 26600 36964
rect 5176 36476 5240 36480
rect 5176 36420 5180 36476
rect 5180 36420 5236 36476
rect 5236 36420 5240 36476
rect 5176 36416 5240 36420
rect 5256 36476 5320 36480
rect 5256 36420 5260 36476
rect 5260 36420 5316 36476
rect 5316 36420 5320 36476
rect 5256 36416 5320 36420
rect 5336 36476 5400 36480
rect 5336 36420 5340 36476
rect 5340 36420 5396 36476
rect 5396 36420 5400 36476
rect 5336 36416 5400 36420
rect 5416 36476 5480 36480
rect 5416 36420 5420 36476
rect 5420 36420 5476 36476
rect 5476 36420 5480 36476
rect 5416 36416 5480 36420
rect 13624 36476 13688 36480
rect 13624 36420 13628 36476
rect 13628 36420 13684 36476
rect 13684 36420 13688 36476
rect 13624 36416 13688 36420
rect 13704 36476 13768 36480
rect 13704 36420 13708 36476
rect 13708 36420 13764 36476
rect 13764 36420 13768 36476
rect 13704 36416 13768 36420
rect 13784 36476 13848 36480
rect 13784 36420 13788 36476
rect 13788 36420 13844 36476
rect 13844 36420 13848 36476
rect 13784 36416 13848 36420
rect 13864 36476 13928 36480
rect 13864 36420 13868 36476
rect 13868 36420 13924 36476
rect 13924 36420 13928 36476
rect 13864 36416 13928 36420
rect 22072 36476 22136 36480
rect 22072 36420 22076 36476
rect 22076 36420 22132 36476
rect 22132 36420 22136 36476
rect 22072 36416 22136 36420
rect 22152 36476 22216 36480
rect 22152 36420 22156 36476
rect 22156 36420 22212 36476
rect 22212 36420 22216 36476
rect 22152 36416 22216 36420
rect 22232 36476 22296 36480
rect 22232 36420 22236 36476
rect 22236 36420 22292 36476
rect 22292 36420 22296 36476
rect 22232 36416 22296 36420
rect 22312 36476 22376 36480
rect 22312 36420 22316 36476
rect 22316 36420 22372 36476
rect 22372 36420 22376 36476
rect 22312 36416 22376 36420
rect 30520 36476 30584 36480
rect 30520 36420 30524 36476
rect 30524 36420 30580 36476
rect 30580 36420 30584 36476
rect 30520 36416 30584 36420
rect 30600 36476 30664 36480
rect 30600 36420 30604 36476
rect 30604 36420 30660 36476
rect 30660 36420 30664 36476
rect 30600 36416 30664 36420
rect 30680 36476 30744 36480
rect 30680 36420 30684 36476
rect 30684 36420 30740 36476
rect 30740 36420 30744 36476
rect 30680 36416 30744 36420
rect 30760 36476 30824 36480
rect 30760 36420 30764 36476
rect 30764 36420 30820 36476
rect 30820 36420 30824 36476
rect 30760 36416 30824 36420
rect 9400 35932 9464 35936
rect 9400 35876 9404 35932
rect 9404 35876 9460 35932
rect 9460 35876 9464 35932
rect 9400 35872 9464 35876
rect 9480 35932 9544 35936
rect 9480 35876 9484 35932
rect 9484 35876 9540 35932
rect 9540 35876 9544 35932
rect 9480 35872 9544 35876
rect 9560 35932 9624 35936
rect 9560 35876 9564 35932
rect 9564 35876 9620 35932
rect 9620 35876 9624 35932
rect 9560 35872 9624 35876
rect 9640 35932 9704 35936
rect 9640 35876 9644 35932
rect 9644 35876 9700 35932
rect 9700 35876 9704 35932
rect 9640 35872 9704 35876
rect 17848 35932 17912 35936
rect 17848 35876 17852 35932
rect 17852 35876 17908 35932
rect 17908 35876 17912 35932
rect 17848 35872 17912 35876
rect 17928 35932 17992 35936
rect 17928 35876 17932 35932
rect 17932 35876 17988 35932
rect 17988 35876 17992 35932
rect 17928 35872 17992 35876
rect 18008 35932 18072 35936
rect 18008 35876 18012 35932
rect 18012 35876 18068 35932
rect 18068 35876 18072 35932
rect 18008 35872 18072 35876
rect 18088 35932 18152 35936
rect 18088 35876 18092 35932
rect 18092 35876 18148 35932
rect 18148 35876 18152 35932
rect 18088 35872 18152 35876
rect 26296 35932 26360 35936
rect 26296 35876 26300 35932
rect 26300 35876 26356 35932
rect 26356 35876 26360 35932
rect 26296 35872 26360 35876
rect 26376 35932 26440 35936
rect 26376 35876 26380 35932
rect 26380 35876 26436 35932
rect 26436 35876 26440 35932
rect 26376 35872 26440 35876
rect 26456 35932 26520 35936
rect 26456 35876 26460 35932
rect 26460 35876 26516 35932
rect 26516 35876 26520 35932
rect 26456 35872 26520 35876
rect 26536 35932 26600 35936
rect 26536 35876 26540 35932
rect 26540 35876 26596 35932
rect 26596 35876 26600 35932
rect 26536 35872 26600 35876
rect 5176 35388 5240 35392
rect 5176 35332 5180 35388
rect 5180 35332 5236 35388
rect 5236 35332 5240 35388
rect 5176 35328 5240 35332
rect 5256 35388 5320 35392
rect 5256 35332 5260 35388
rect 5260 35332 5316 35388
rect 5316 35332 5320 35388
rect 5256 35328 5320 35332
rect 5336 35388 5400 35392
rect 5336 35332 5340 35388
rect 5340 35332 5396 35388
rect 5396 35332 5400 35388
rect 5336 35328 5400 35332
rect 5416 35388 5480 35392
rect 5416 35332 5420 35388
rect 5420 35332 5476 35388
rect 5476 35332 5480 35388
rect 5416 35328 5480 35332
rect 13624 35388 13688 35392
rect 13624 35332 13628 35388
rect 13628 35332 13684 35388
rect 13684 35332 13688 35388
rect 13624 35328 13688 35332
rect 13704 35388 13768 35392
rect 13704 35332 13708 35388
rect 13708 35332 13764 35388
rect 13764 35332 13768 35388
rect 13704 35328 13768 35332
rect 13784 35388 13848 35392
rect 13784 35332 13788 35388
rect 13788 35332 13844 35388
rect 13844 35332 13848 35388
rect 13784 35328 13848 35332
rect 13864 35388 13928 35392
rect 13864 35332 13868 35388
rect 13868 35332 13924 35388
rect 13924 35332 13928 35388
rect 13864 35328 13928 35332
rect 22072 35388 22136 35392
rect 22072 35332 22076 35388
rect 22076 35332 22132 35388
rect 22132 35332 22136 35388
rect 22072 35328 22136 35332
rect 22152 35388 22216 35392
rect 22152 35332 22156 35388
rect 22156 35332 22212 35388
rect 22212 35332 22216 35388
rect 22152 35328 22216 35332
rect 22232 35388 22296 35392
rect 22232 35332 22236 35388
rect 22236 35332 22292 35388
rect 22292 35332 22296 35388
rect 22232 35328 22296 35332
rect 22312 35388 22376 35392
rect 22312 35332 22316 35388
rect 22316 35332 22372 35388
rect 22372 35332 22376 35388
rect 22312 35328 22376 35332
rect 30520 35388 30584 35392
rect 30520 35332 30524 35388
rect 30524 35332 30580 35388
rect 30580 35332 30584 35388
rect 30520 35328 30584 35332
rect 30600 35388 30664 35392
rect 30600 35332 30604 35388
rect 30604 35332 30660 35388
rect 30660 35332 30664 35388
rect 30600 35328 30664 35332
rect 30680 35388 30744 35392
rect 30680 35332 30684 35388
rect 30684 35332 30740 35388
rect 30740 35332 30744 35388
rect 30680 35328 30744 35332
rect 30760 35388 30824 35392
rect 30760 35332 30764 35388
rect 30764 35332 30820 35388
rect 30820 35332 30824 35388
rect 30760 35328 30824 35332
rect 9400 34844 9464 34848
rect 9400 34788 9404 34844
rect 9404 34788 9460 34844
rect 9460 34788 9464 34844
rect 9400 34784 9464 34788
rect 9480 34844 9544 34848
rect 9480 34788 9484 34844
rect 9484 34788 9540 34844
rect 9540 34788 9544 34844
rect 9480 34784 9544 34788
rect 9560 34844 9624 34848
rect 9560 34788 9564 34844
rect 9564 34788 9620 34844
rect 9620 34788 9624 34844
rect 9560 34784 9624 34788
rect 9640 34844 9704 34848
rect 9640 34788 9644 34844
rect 9644 34788 9700 34844
rect 9700 34788 9704 34844
rect 9640 34784 9704 34788
rect 17848 34844 17912 34848
rect 17848 34788 17852 34844
rect 17852 34788 17908 34844
rect 17908 34788 17912 34844
rect 17848 34784 17912 34788
rect 17928 34844 17992 34848
rect 17928 34788 17932 34844
rect 17932 34788 17988 34844
rect 17988 34788 17992 34844
rect 17928 34784 17992 34788
rect 18008 34844 18072 34848
rect 18008 34788 18012 34844
rect 18012 34788 18068 34844
rect 18068 34788 18072 34844
rect 18008 34784 18072 34788
rect 18088 34844 18152 34848
rect 18088 34788 18092 34844
rect 18092 34788 18148 34844
rect 18148 34788 18152 34844
rect 18088 34784 18152 34788
rect 26296 34844 26360 34848
rect 26296 34788 26300 34844
rect 26300 34788 26356 34844
rect 26356 34788 26360 34844
rect 26296 34784 26360 34788
rect 26376 34844 26440 34848
rect 26376 34788 26380 34844
rect 26380 34788 26436 34844
rect 26436 34788 26440 34844
rect 26376 34784 26440 34788
rect 26456 34844 26520 34848
rect 26456 34788 26460 34844
rect 26460 34788 26516 34844
rect 26516 34788 26520 34844
rect 26456 34784 26520 34788
rect 26536 34844 26600 34848
rect 26536 34788 26540 34844
rect 26540 34788 26596 34844
rect 26596 34788 26600 34844
rect 26536 34784 26600 34788
rect 5176 34300 5240 34304
rect 5176 34244 5180 34300
rect 5180 34244 5236 34300
rect 5236 34244 5240 34300
rect 5176 34240 5240 34244
rect 5256 34300 5320 34304
rect 5256 34244 5260 34300
rect 5260 34244 5316 34300
rect 5316 34244 5320 34300
rect 5256 34240 5320 34244
rect 5336 34300 5400 34304
rect 5336 34244 5340 34300
rect 5340 34244 5396 34300
rect 5396 34244 5400 34300
rect 5336 34240 5400 34244
rect 5416 34300 5480 34304
rect 5416 34244 5420 34300
rect 5420 34244 5476 34300
rect 5476 34244 5480 34300
rect 5416 34240 5480 34244
rect 13624 34300 13688 34304
rect 13624 34244 13628 34300
rect 13628 34244 13684 34300
rect 13684 34244 13688 34300
rect 13624 34240 13688 34244
rect 13704 34300 13768 34304
rect 13704 34244 13708 34300
rect 13708 34244 13764 34300
rect 13764 34244 13768 34300
rect 13704 34240 13768 34244
rect 13784 34300 13848 34304
rect 13784 34244 13788 34300
rect 13788 34244 13844 34300
rect 13844 34244 13848 34300
rect 13784 34240 13848 34244
rect 13864 34300 13928 34304
rect 13864 34244 13868 34300
rect 13868 34244 13924 34300
rect 13924 34244 13928 34300
rect 13864 34240 13928 34244
rect 22072 34300 22136 34304
rect 22072 34244 22076 34300
rect 22076 34244 22132 34300
rect 22132 34244 22136 34300
rect 22072 34240 22136 34244
rect 22152 34300 22216 34304
rect 22152 34244 22156 34300
rect 22156 34244 22212 34300
rect 22212 34244 22216 34300
rect 22152 34240 22216 34244
rect 22232 34300 22296 34304
rect 22232 34244 22236 34300
rect 22236 34244 22292 34300
rect 22292 34244 22296 34300
rect 22232 34240 22296 34244
rect 22312 34300 22376 34304
rect 22312 34244 22316 34300
rect 22316 34244 22372 34300
rect 22372 34244 22376 34300
rect 22312 34240 22376 34244
rect 30520 34300 30584 34304
rect 30520 34244 30524 34300
rect 30524 34244 30580 34300
rect 30580 34244 30584 34300
rect 30520 34240 30584 34244
rect 30600 34300 30664 34304
rect 30600 34244 30604 34300
rect 30604 34244 30660 34300
rect 30660 34244 30664 34300
rect 30600 34240 30664 34244
rect 30680 34300 30744 34304
rect 30680 34244 30684 34300
rect 30684 34244 30740 34300
rect 30740 34244 30744 34300
rect 30680 34240 30744 34244
rect 30760 34300 30824 34304
rect 30760 34244 30764 34300
rect 30764 34244 30820 34300
rect 30820 34244 30824 34300
rect 30760 34240 30824 34244
rect 9400 33756 9464 33760
rect 9400 33700 9404 33756
rect 9404 33700 9460 33756
rect 9460 33700 9464 33756
rect 9400 33696 9464 33700
rect 9480 33756 9544 33760
rect 9480 33700 9484 33756
rect 9484 33700 9540 33756
rect 9540 33700 9544 33756
rect 9480 33696 9544 33700
rect 9560 33756 9624 33760
rect 9560 33700 9564 33756
rect 9564 33700 9620 33756
rect 9620 33700 9624 33756
rect 9560 33696 9624 33700
rect 9640 33756 9704 33760
rect 9640 33700 9644 33756
rect 9644 33700 9700 33756
rect 9700 33700 9704 33756
rect 9640 33696 9704 33700
rect 17848 33756 17912 33760
rect 17848 33700 17852 33756
rect 17852 33700 17908 33756
rect 17908 33700 17912 33756
rect 17848 33696 17912 33700
rect 17928 33756 17992 33760
rect 17928 33700 17932 33756
rect 17932 33700 17988 33756
rect 17988 33700 17992 33756
rect 17928 33696 17992 33700
rect 18008 33756 18072 33760
rect 18008 33700 18012 33756
rect 18012 33700 18068 33756
rect 18068 33700 18072 33756
rect 18008 33696 18072 33700
rect 18088 33756 18152 33760
rect 18088 33700 18092 33756
rect 18092 33700 18148 33756
rect 18148 33700 18152 33756
rect 18088 33696 18152 33700
rect 26296 33756 26360 33760
rect 26296 33700 26300 33756
rect 26300 33700 26356 33756
rect 26356 33700 26360 33756
rect 26296 33696 26360 33700
rect 26376 33756 26440 33760
rect 26376 33700 26380 33756
rect 26380 33700 26436 33756
rect 26436 33700 26440 33756
rect 26376 33696 26440 33700
rect 26456 33756 26520 33760
rect 26456 33700 26460 33756
rect 26460 33700 26516 33756
rect 26516 33700 26520 33756
rect 26456 33696 26520 33700
rect 26536 33756 26600 33760
rect 26536 33700 26540 33756
rect 26540 33700 26596 33756
rect 26596 33700 26600 33756
rect 26536 33696 26600 33700
rect 5176 33212 5240 33216
rect 5176 33156 5180 33212
rect 5180 33156 5236 33212
rect 5236 33156 5240 33212
rect 5176 33152 5240 33156
rect 5256 33212 5320 33216
rect 5256 33156 5260 33212
rect 5260 33156 5316 33212
rect 5316 33156 5320 33212
rect 5256 33152 5320 33156
rect 5336 33212 5400 33216
rect 5336 33156 5340 33212
rect 5340 33156 5396 33212
rect 5396 33156 5400 33212
rect 5336 33152 5400 33156
rect 5416 33212 5480 33216
rect 5416 33156 5420 33212
rect 5420 33156 5476 33212
rect 5476 33156 5480 33212
rect 5416 33152 5480 33156
rect 13624 33212 13688 33216
rect 13624 33156 13628 33212
rect 13628 33156 13684 33212
rect 13684 33156 13688 33212
rect 13624 33152 13688 33156
rect 13704 33212 13768 33216
rect 13704 33156 13708 33212
rect 13708 33156 13764 33212
rect 13764 33156 13768 33212
rect 13704 33152 13768 33156
rect 13784 33212 13848 33216
rect 13784 33156 13788 33212
rect 13788 33156 13844 33212
rect 13844 33156 13848 33212
rect 13784 33152 13848 33156
rect 13864 33212 13928 33216
rect 13864 33156 13868 33212
rect 13868 33156 13924 33212
rect 13924 33156 13928 33212
rect 13864 33152 13928 33156
rect 22072 33212 22136 33216
rect 22072 33156 22076 33212
rect 22076 33156 22132 33212
rect 22132 33156 22136 33212
rect 22072 33152 22136 33156
rect 22152 33212 22216 33216
rect 22152 33156 22156 33212
rect 22156 33156 22212 33212
rect 22212 33156 22216 33212
rect 22152 33152 22216 33156
rect 22232 33212 22296 33216
rect 22232 33156 22236 33212
rect 22236 33156 22292 33212
rect 22292 33156 22296 33212
rect 22232 33152 22296 33156
rect 22312 33212 22376 33216
rect 22312 33156 22316 33212
rect 22316 33156 22372 33212
rect 22372 33156 22376 33212
rect 22312 33152 22376 33156
rect 30520 33212 30584 33216
rect 30520 33156 30524 33212
rect 30524 33156 30580 33212
rect 30580 33156 30584 33212
rect 30520 33152 30584 33156
rect 30600 33212 30664 33216
rect 30600 33156 30604 33212
rect 30604 33156 30660 33212
rect 30660 33156 30664 33212
rect 30600 33152 30664 33156
rect 30680 33212 30744 33216
rect 30680 33156 30684 33212
rect 30684 33156 30740 33212
rect 30740 33156 30744 33212
rect 30680 33152 30744 33156
rect 30760 33212 30824 33216
rect 30760 33156 30764 33212
rect 30764 33156 30820 33212
rect 30820 33156 30824 33212
rect 30760 33152 30824 33156
rect 9400 32668 9464 32672
rect 9400 32612 9404 32668
rect 9404 32612 9460 32668
rect 9460 32612 9464 32668
rect 9400 32608 9464 32612
rect 9480 32668 9544 32672
rect 9480 32612 9484 32668
rect 9484 32612 9540 32668
rect 9540 32612 9544 32668
rect 9480 32608 9544 32612
rect 9560 32668 9624 32672
rect 9560 32612 9564 32668
rect 9564 32612 9620 32668
rect 9620 32612 9624 32668
rect 9560 32608 9624 32612
rect 9640 32668 9704 32672
rect 9640 32612 9644 32668
rect 9644 32612 9700 32668
rect 9700 32612 9704 32668
rect 9640 32608 9704 32612
rect 17848 32668 17912 32672
rect 17848 32612 17852 32668
rect 17852 32612 17908 32668
rect 17908 32612 17912 32668
rect 17848 32608 17912 32612
rect 17928 32668 17992 32672
rect 17928 32612 17932 32668
rect 17932 32612 17988 32668
rect 17988 32612 17992 32668
rect 17928 32608 17992 32612
rect 18008 32668 18072 32672
rect 18008 32612 18012 32668
rect 18012 32612 18068 32668
rect 18068 32612 18072 32668
rect 18008 32608 18072 32612
rect 18088 32668 18152 32672
rect 18088 32612 18092 32668
rect 18092 32612 18148 32668
rect 18148 32612 18152 32668
rect 18088 32608 18152 32612
rect 26296 32668 26360 32672
rect 26296 32612 26300 32668
rect 26300 32612 26356 32668
rect 26356 32612 26360 32668
rect 26296 32608 26360 32612
rect 26376 32668 26440 32672
rect 26376 32612 26380 32668
rect 26380 32612 26436 32668
rect 26436 32612 26440 32668
rect 26376 32608 26440 32612
rect 26456 32668 26520 32672
rect 26456 32612 26460 32668
rect 26460 32612 26516 32668
rect 26516 32612 26520 32668
rect 26456 32608 26520 32612
rect 26536 32668 26600 32672
rect 26536 32612 26540 32668
rect 26540 32612 26596 32668
rect 26596 32612 26600 32668
rect 26536 32608 26600 32612
rect 5176 32124 5240 32128
rect 5176 32068 5180 32124
rect 5180 32068 5236 32124
rect 5236 32068 5240 32124
rect 5176 32064 5240 32068
rect 5256 32124 5320 32128
rect 5256 32068 5260 32124
rect 5260 32068 5316 32124
rect 5316 32068 5320 32124
rect 5256 32064 5320 32068
rect 5336 32124 5400 32128
rect 5336 32068 5340 32124
rect 5340 32068 5396 32124
rect 5396 32068 5400 32124
rect 5336 32064 5400 32068
rect 5416 32124 5480 32128
rect 5416 32068 5420 32124
rect 5420 32068 5476 32124
rect 5476 32068 5480 32124
rect 5416 32064 5480 32068
rect 13624 32124 13688 32128
rect 13624 32068 13628 32124
rect 13628 32068 13684 32124
rect 13684 32068 13688 32124
rect 13624 32064 13688 32068
rect 13704 32124 13768 32128
rect 13704 32068 13708 32124
rect 13708 32068 13764 32124
rect 13764 32068 13768 32124
rect 13704 32064 13768 32068
rect 13784 32124 13848 32128
rect 13784 32068 13788 32124
rect 13788 32068 13844 32124
rect 13844 32068 13848 32124
rect 13784 32064 13848 32068
rect 13864 32124 13928 32128
rect 13864 32068 13868 32124
rect 13868 32068 13924 32124
rect 13924 32068 13928 32124
rect 13864 32064 13928 32068
rect 22072 32124 22136 32128
rect 22072 32068 22076 32124
rect 22076 32068 22132 32124
rect 22132 32068 22136 32124
rect 22072 32064 22136 32068
rect 22152 32124 22216 32128
rect 22152 32068 22156 32124
rect 22156 32068 22212 32124
rect 22212 32068 22216 32124
rect 22152 32064 22216 32068
rect 22232 32124 22296 32128
rect 22232 32068 22236 32124
rect 22236 32068 22292 32124
rect 22292 32068 22296 32124
rect 22232 32064 22296 32068
rect 22312 32124 22376 32128
rect 22312 32068 22316 32124
rect 22316 32068 22372 32124
rect 22372 32068 22376 32124
rect 22312 32064 22376 32068
rect 30520 32124 30584 32128
rect 30520 32068 30524 32124
rect 30524 32068 30580 32124
rect 30580 32068 30584 32124
rect 30520 32064 30584 32068
rect 30600 32124 30664 32128
rect 30600 32068 30604 32124
rect 30604 32068 30660 32124
rect 30660 32068 30664 32124
rect 30600 32064 30664 32068
rect 30680 32124 30744 32128
rect 30680 32068 30684 32124
rect 30684 32068 30740 32124
rect 30740 32068 30744 32124
rect 30680 32064 30744 32068
rect 30760 32124 30824 32128
rect 30760 32068 30764 32124
rect 30764 32068 30820 32124
rect 30820 32068 30824 32124
rect 30760 32064 30824 32068
rect 9400 31580 9464 31584
rect 9400 31524 9404 31580
rect 9404 31524 9460 31580
rect 9460 31524 9464 31580
rect 9400 31520 9464 31524
rect 9480 31580 9544 31584
rect 9480 31524 9484 31580
rect 9484 31524 9540 31580
rect 9540 31524 9544 31580
rect 9480 31520 9544 31524
rect 9560 31580 9624 31584
rect 9560 31524 9564 31580
rect 9564 31524 9620 31580
rect 9620 31524 9624 31580
rect 9560 31520 9624 31524
rect 9640 31580 9704 31584
rect 9640 31524 9644 31580
rect 9644 31524 9700 31580
rect 9700 31524 9704 31580
rect 9640 31520 9704 31524
rect 17848 31580 17912 31584
rect 17848 31524 17852 31580
rect 17852 31524 17908 31580
rect 17908 31524 17912 31580
rect 17848 31520 17912 31524
rect 17928 31580 17992 31584
rect 17928 31524 17932 31580
rect 17932 31524 17988 31580
rect 17988 31524 17992 31580
rect 17928 31520 17992 31524
rect 18008 31580 18072 31584
rect 18008 31524 18012 31580
rect 18012 31524 18068 31580
rect 18068 31524 18072 31580
rect 18008 31520 18072 31524
rect 18088 31580 18152 31584
rect 18088 31524 18092 31580
rect 18092 31524 18148 31580
rect 18148 31524 18152 31580
rect 18088 31520 18152 31524
rect 26296 31580 26360 31584
rect 26296 31524 26300 31580
rect 26300 31524 26356 31580
rect 26356 31524 26360 31580
rect 26296 31520 26360 31524
rect 26376 31580 26440 31584
rect 26376 31524 26380 31580
rect 26380 31524 26436 31580
rect 26436 31524 26440 31580
rect 26376 31520 26440 31524
rect 26456 31580 26520 31584
rect 26456 31524 26460 31580
rect 26460 31524 26516 31580
rect 26516 31524 26520 31580
rect 26456 31520 26520 31524
rect 26536 31580 26600 31584
rect 26536 31524 26540 31580
rect 26540 31524 26596 31580
rect 26596 31524 26600 31580
rect 26536 31520 26600 31524
rect 5176 31036 5240 31040
rect 5176 30980 5180 31036
rect 5180 30980 5236 31036
rect 5236 30980 5240 31036
rect 5176 30976 5240 30980
rect 5256 31036 5320 31040
rect 5256 30980 5260 31036
rect 5260 30980 5316 31036
rect 5316 30980 5320 31036
rect 5256 30976 5320 30980
rect 5336 31036 5400 31040
rect 5336 30980 5340 31036
rect 5340 30980 5396 31036
rect 5396 30980 5400 31036
rect 5336 30976 5400 30980
rect 5416 31036 5480 31040
rect 5416 30980 5420 31036
rect 5420 30980 5476 31036
rect 5476 30980 5480 31036
rect 5416 30976 5480 30980
rect 13624 31036 13688 31040
rect 13624 30980 13628 31036
rect 13628 30980 13684 31036
rect 13684 30980 13688 31036
rect 13624 30976 13688 30980
rect 13704 31036 13768 31040
rect 13704 30980 13708 31036
rect 13708 30980 13764 31036
rect 13764 30980 13768 31036
rect 13704 30976 13768 30980
rect 13784 31036 13848 31040
rect 13784 30980 13788 31036
rect 13788 30980 13844 31036
rect 13844 30980 13848 31036
rect 13784 30976 13848 30980
rect 13864 31036 13928 31040
rect 13864 30980 13868 31036
rect 13868 30980 13924 31036
rect 13924 30980 13928 31036
rect 13864 30976 13928 30980
rect 22072 31036 22136 31040
rect 22072 30980 22076 31036
rect 22076 30980 22132 31036
rect 22132 30980 22136 31036
rect 22072 30976 22136 30980
rect 22152 31036 22216 31040
rect 22152 30980 22156 31036
rect 22156 30980 22212 31036
rect 22212 30980 22216 31036
rect 22152 30976 22216 30980
rect 22232 31036 22296 31040
rect 22232 30980 22236 31036
rect 22236 30980 22292 31036
rect 22292 30980 22296 31036
rect 22232 30976 22296 30980
rect 22312 31036 22376 31040
rect 22312 30980 22316 31036
rect 22316 30980 22372 31036
rect 22372 30980 22376 31036
rect 22312 30976 22376 30980
rect 30520 31036 30584 31040
rect 30520 30980 30524 31036
rect 30524 30980 30580 31036
rect 30580 30980 30584 31036
rect 30520 30976 30584 30980
rect 30600 31036 30664 31040
rect 30600 30980 30604 31036
rect 30604 30980 30660 31036
rect 30660 30980 30664 31036
rect 30600 30976 30664 30980
rect 30680 31036 30744 31040
rect 30680 30980 30684 31036
rect 30684 30980 30740 31036
rect 30740 30980 30744 31036
rect 30680 30976 30744 30980
rect 30760 31036 30824 31040
rect 30760 30980 30764 31036
rect 30764 30980 30820 31036
rect 30820 30980 30824 31036
rect 30760 30976 30824 30980
rect 9400 30492 9464 30496
rect 9400 30436 9404 30492
rect 9404 30436 9460 30492
rect 9460 30436 9464 30492
rect 9400 30432 9464 30436
rect 9480 30492 9544 30496
rect 9480 30436 9484 30492
rect 9484 30436 9540 30492
rect 9540 30436 9544 30492
rect 9480 30432 9544 30436
rect 9560 30492 9624 30496
rect 9560 30436 9564 30492
rect 9564 30436 9620 30492
rect 9620 30436 9624 30492
rect 9560 30432 9624 30436
rect 9640 30492 9704 30496
rect 9640 30436 9644 30492
rect 9644 30436 9700 30492
rect 9700 30436 9704 30492
rect 9640 30432 9704 30436
rect 17848 30492 17912 30496
rect 17848 30436 17852 30492
rect 17852 30436 17908 30492
rect 17908 30436 17912 30492
rect 17848 30432 17912 30436
rect 17928 30492 17992 30496
rect 17928 30436 17932 30492
rect 17932 30436 17988 30492
rect 17988 30436 17992 30492
rect 17928 30432 17992 30436
rect 18008 30492 18072 30496
rect 18008 30436 18012 30492
rect 18012 30436 18068 30492
rect 18068 30436 18072 30492
rect 18008 30432 18072 30436
rect 18088 30492 18152 30496
rect 18088 30436 18092 30492
rect 18092 30436 18148 30492
rect 18148 30436 18152 30492
rect 18088 30432 18152 30436
rect 26296 30492 26360 30496
rect 26296 30436 26300 30492
rect 26300 30436 26356 30492
rect 26356 30436 26360 30492
rect 26296 30432 26360 30436
rect 26376 30492 26440 30496
rect 26376 30436 26380 30492
rect 26380 30436 26436 30492
rect 26436 30436 26440 30492
rect 26376 30432 26440 30436
rect 26456 30492 26520 30496
rect 26456 30436 26460 30492
rect 26460 30436 26516 30492
rect 26516 30436 26520 30492
rect 26456 30432 26520 30436
rect 26536 30492 26600 30496
rect 26536 30436 26540 30492
rect 26540 30436 26596 30492
rect 26596 30436 26600 30492
rect 26536 30432 26600 30436
rect 5176 29948 5240 29952
rect 5176 29892 5180 29948
rect 5180 29892 5236 29948
rect 5236 29892 5240 29948
rect 5176 29888 5240 29892
rect 5256 29948 5320 29952
rect 5256 29892 5260 29948
rect 5260 29892 5316 29948
rect 5316 29892 5320 29948
rect 5256 29888 5320 29892
rect 5336 29948 5400 29952
rect 5336 29892 5340 29948
rect 5340 29892 5396 29948
rect 5396 29892 5400 29948
rect 5336 29888 5400 29892
rect 5416 29948 5480 29952
rect 5416 29892 5420 29948
rect 5420 29892 5476 29948
rect 5476 29892 5480 29948
rect 5416 29888 5480 29892
rect 13624 29948 13688 29952
rect 13624 29892 13628 29948
rect 13628 29892 13684 29948
rect 13684 29892 13688 29948
rect 13624 29888 13688 29892
rect 13704 29948 13768 29952
rect 13704 29892 13708 29948
rect 13708 29892 13764 29948
rect 13764 29892 13768 29948
rect 13704 29888 13768 29892
rect 13784 29948 13848 29952
rect 13784 29892 13788 29948
rect 13788 29892 13844 29948
rect 13844 29892 13848 29948
rect 13784 29888 13848 29892
rect 13864 29948 13928 29952
rect 13864 29892 13868 29948
rect 13868 29892 13924 29948
rect 13924 29892 13928 29948
rect 13864 29888 13928 29892
rect 22072 29948 22136 29952
rect 22072 29892 22076 29948
rect 22076 29892 22132 29948
rect 22132 29892 22136 29948
rect 22072 29888 22136 29892
rect 22152 29948 22216 29952
rect 22152 29892 22156 29948
rect 22156 29892 22212 29948
rect 22212 29892 22216 29948
rect 22152 29888 22216 29892
rect 22232 29948 22296 29952
rect 22232 29892 22236 29948
rect 22236 29892 22292 29948
rect 22292 29892 22296 29948
rect 22232 29888 22296 29892
rect 22312 29948 22376 29952
rect 22312 29892 22316 29948
rect 22316 29892 22372 29948
rect 22372 29892 22376 29948
rect 22312 29888 22376 29892
rect 30520 29948 30584 29952
rect 30520 29892 30524 29948
rect 30524 29892 30580 29948
rect 30580 29892 30584 29948
rect 30520 29888 30584 29892
rect 30600 29948 30664 29952
rect 30600 29892 30604 29948
rect 30604 29892 30660 29948
rect 30660 29892 30664 29948
rect 30600 29888 30664 29892
rect 30680 29948 30744 29952
rect 30680 29892 30684 29948
rect 30684 29892 30740 29948
rect 30740 29892 30744 29948
rect 30680 29888 30744 29892
rect 30760 29948 30824 29952
rect 30760 29892 30764 29948
rect 30764 29892 30820 29948
rect 30820 29892 30824 29948
rect 30760 29888 30824 29892
rect 9400 29404 9464 29408
rect 9400 29348 9404 29404
rect 9404 29348 9460 29404
rect 9460 29348 9464 29404
rect 9400 29344 9464 29348
rect 9480 29404 9544 29408
rect 9480 29348 9484 29404
rect 9484 29348 9540 29404
rect 9540 29348 9544 29404
rect 9480 29344 9544 29348
rect 9560 29404 9624 29408
rect 9560 29348 9564 29404
rect 9564 29348 9620 29404
rect 9620 29348 9624 29404
rect 9560 29344 9624 29348
rect 9640 29404 9704 29408
rect 9640 29348 9644 29404
rect 9644 29348 9700 29404
rect 9700 29348 9704 29404
rect 9640 29344 9704 29348
rect 17848 29404 17912 29408
rect 17848 29348 17852 29404
rect 17852 29348 17908 29404
rect 17908 29348 17912 29404
rect 17848 29344 17912 29348
rect 17928 29404 17992 29408
rect 17928 29348 17932 29404
rect 17932 29348 17988 29404
rect 17988 29348 17992 29404
rect 17928 29344 17992 29348
rect 18008 29404 18072 29408
rect 18008 29348 18012 29404
rect 18012 29348 18068 29404
rect 18068 29348 18072 29404
rect 18008 29344 18072 29348
rect 18088 29404 18152 29408
rect 18088 29348 18092 29404
rect 18092 29348 18148 29404
rect 18148 29348 18152 29404
rect 18088 29344 18152 29348
rect 26296 29404 26360 29408
rect 26296 29348 26300 29404
rect 26300 29348 26356 29404
rect 26356 29348 26360 29404
rect 26296 29344 26360 29348
rect 26376 29404 26440 29408
rect 26376 29348 26380 29404
rect 26380 29348 26436 29404
rect 26436 29348 26440 29404
rect 26376 29344 26440 29348
rect 26456 29404 26520 29408
rect 26456 29348 26460 29404
rect 26460 29348 26516 29404
rect 26516 29348 26520 29404
rect 26456 29344 26520 29348
rect 26536 29404 26600 29408
rect 26536 29348 26540 29404
rect 26540 29348 26596 29404
rect 26596 29348 26600 29404
rect 26536 29344 26600 29348
rect 5176 28860 5240 28864
rect 5176 28804 5180 28860
rect 5180 28804 5236 28860
rect 5236 28804 5240 28860
rect 5176 28800 5240 28804
rect 5256 28860 5320 28864
rect 5256 28804 5260 28860
rect 5260 28804 5316 28860
rect 5316 28804 5320 28860
rect 5256 28800 5320 28804
rect 5336 28860 5400 28864
rect 5336 28804 5340 28860
rect 5340 28804 5396 28860
rect 5396 28804 5400 28860
rect 5336 28800 5400 28804
rect 5416 28860 5480 28864
rect 5416 28804 5420 28860
rect 5420 28804 5476 28860
rect 5476 28804 5480 28860
rect 5416 28800 5480 28804
rect 13624 28860 13688 28864
rect 13624 28804 13628 28860
rect 13628 28804 13684 28860
rect 13684 28804 13688 28860
rect 13624 28800 13688 28804
rect 13704 28860 13768 28864
rect 13704 28804 13708 28860
rect 13708 28804 13764 28860
rect 13764 28804 13768 28860
rect 13704 28800 13768 28804
rect 13784 28860 13848 28864
rect 13784 28804 13788 28860
rect 13788 28804 13844 28860
rect 13844 28804 13848 28860
rect 13784 28800 13848 28804
rect 13864 28860 13928 28864
rect 13864 28804 13868 28860
rect 13868 28804 13924 28860
rect 13924 28804 13928 28860
rect 13864 28800 13928 28804
rect 22072 28860 22136 28864
rect 22072 28804 22076 28860
rect 22076 28804 22132 28860
rect 22132 28804 22136 28860
rect 22072 28800 22136 28804
rect 22152 28860 22216 28864
rect 22152 28804 22156 28860
rect 22156 28804 22212 28860
rect 22212 28804 22216 28860
rect 22152 28800 22216 28804
rect 22232 28860 22296 28864
rect 22232 28804 22236 28860
rect 22236 28804 22292 28860
rect 22292 28804 22296 28860
rect 22232 28800 22296 28804
rect 22312 28860 22376 28864
rect 22312 28804 22316 28860
rect 22316 28804 22372 28860
rect 22372 28804 22376 28860
rect 22312 28800 22376 28804
rect 30520 28860 30584 28864
rect 30520 28804 30524 28860
rect 30524 28804 30580 28860
rect 30580 28804 30584 28860
rect 30520 28800 30584 28804
rect 30600 28860 30664 28864
rect 30600 28804 30604 28860
rect 30604 28804 30660 28860
rect 30660 28804 30664 28860
rect 30600 28800 30664 28804
rect 30680 28860 30744 28864
rect 30680 28804 30684 28860
rect 30684 28804 30740 28860
rect 30740 28804 30744 28860
rect 30680 28800 30744 28804
rect 30760 28860 30824 28864
rect 30760 28804 30764 28860
rect 30764 28804 30820 28860
rect 30820 28804 30824 28860
rect 30760 28800 30824 28804
rect 9400 28316 9464 28320
rect 9400 28260 9404 28316
rect 9404 28260 9460 28316
rect 9460 28260 9464 28316
rect 9400 28256 9464 28260
rect 9480 28316 9544 28320
rect 9480 28260 9484 28316
rect 9484 28260 9540 28316
rect 9540 28260 9544 28316
rect 9480 28256 9544 28260
rect 9560 28316 9624 28320
rect 9560 28260 9564 28316
rect 9564 28260 9620 28316
rect 9620 28260 9624 28316
rect 9560 28256 9624 28260
rect 9640 28316 9704 28320
rect 9640 28260 9644 28316
rect 9644 28260 9700 28316
rect 9700 28260 9704 28316
rect 9640 28256 9704 28260
rect 17848 28316 17912 28320
rect 17848 28260 17852 28316
rect 17852 28260 17908 28316
rect 17908 28260 17912 28316
rect 17848 28256 17912 28260
rect 17928 28316 17992 28320
rect 17928 28260 17932 28316
rect 17932 28260 17988 28316
rect 17988 28260 17992 28316
rect 17928 28256 17992 28260
rect 18008 28316 18072 28320
rect 18008 28260 18012 28316
rect 18012 28260 18068 28316
rect 18068 28260 18072 28316
rect 18008 28256 18072 28260
rect 18088 28316 18152 28320
rect 18088 28260 18092 28316
rect 18092 28260 18148 28316
rect 18148 28260 18152 28316
rect 18088 28256 18152 28260
rect 26296 28316 26360 28320
rect 26296 28260 26300 28316
rect 26300 28260 26356 28316
rect 26356 28260 26360 28316
rect 26296 28256 26360 28260
rect 26376 28316 26440 28320
rect 26376 28260 26380 28316
rect 26380 28260 26436 28316
rect 26436 28260 26440 28316
rect 26376 28256 26440 28260
rect 26456 28316 26520 28320
rect 26456 28260 26460 28316
rect 26460 28260 26516 28316
rect 26516 28260 26520 28316
rect 26456 28256 26520 28260
rect 26536 28316 26600 28320
rect 26536 28260 26540 28316
rect 26540 28260 26596 28316
rect 26596 28260 26600 28316
rect 26536 28256 26600 28260
rect 5176 27772 5240 27776
rect 5176 27716 5180 27772
rect 5180 27716 5236 27772
rect 5236 27716 5240 27772
rect 5176 27712 5240 27716
rect 5256 27772 5320 27776
rect 5256 27716 5260 27772
rect 5260 27716 5316 27772
rect 5316 27716 5320 27772
rect 5256 27712 5320 27716
rect 5336 27772 5400 27776
rect 5336 27716 5340 27772
rect 5340 27716 5396 27772
rect 5396 27716 5400 27772
rect 5336 27712 5400 27716
rect 5416 27772 5480 27776
rect 5416 27716 5420 27772
rect 5420 27716 5476 27772
rect 5476 27716 5480 27772
rect 5416 27712 5480 27716
rect 13624 27772 13688 27776
rect 13624 27716 13628 27772
rect 13628 27716 13684 27772
rect 13684 27716 13688 27772
rect 13624 27712 13688 27716
rect 13704 27772 13768 27776
rect 13704 27716 13708 27772
rect 13708 27716 13764 27772
rect 13764 27716 13768 27772
rect 13704 27712 13768 27716
rect 13784 27772 13848 27776
rect 13784 27716 13788 27772
rect 13788 27716 13844 27772
rect 13844 27716 13848 27772
rect 13784 27712 13848 27716
rect 13864 27772 13928 27776
rect 13864 27716 13868 27772
rect 13868 27716 13924 27772
rect 13924 27716 13928 27772
rect 13864 27712 13928 27716
rect 22072 27772 22136 27776
rect 22072 27716 22076 27772
rect 22076 27716 22132 27772
rect 22132 27716 22136 27772
rect 22072 27712 22136 27716
rect 22152 27772 22216 27776
rect 22152 27716 22156 27772
rect 22156 27716 22212 27772
rect 22212 27716 22216 27772
rect 22152 27712 22216 27716
rect 22232 27772 22296 27776
rect 22232 27716 22236 27772
rect 22236 27716 22292 27772
rect 22292 27716 22296 27772
rect 22232 27712 22296 27716
rect 22312 27772 22376 27776
rect 22312 27716 22316 27772
rect 22316 27716 22372 27772
rect 22372 27716 22376 27772
rect 22312 27712 22376 27716
rect 30520 27772 30584 27776
rect 30520 27716 30524 27772
rect 30524 27716 30580 27772
rect 30580 27716 30584 27772
rect 30520 27712 30584 27716
rect 30600 27772 30664 27776
rect 30600 27716 30604 27772
rect 30604 27716 30660 27772
rect 30660 27716 30664 27772
rect 30600 27712 30664 27716
rect 30680 27772 30744 27776
rect 30680 27716 30684 27772
rect 30684 27716 30740 27772
rect 30740 27716 30744 27772
rect 30680 27712 30744 27716
rect 30760 27772 30824 27776
rect 30760 27716 30764 27772
rect 30764 27716 30820 27772
rect 30820 27716 30824 27772
rect 30760 27712 30824 27716
rect 9400 27228 9464 27232
rect 9400 27172 9404 27228
rect 9404 27172 9460 27228
rect 9460 27172 9464 27228
rect 9400 27168 9464 27172
rect 9480 27228 9544 27232
rect 9480 27172 9484 27228
rect 9484 27172 9540 27228
rect 9540 27172 9544 27228
rect 9480 27168 9544 27172
rect 9560 27228 9624 27232
rect 9560 27172 9564 27228
rect 9564 27172 9620 27228
rect 9620 27172 9624 27228
rect 9560 27168 9624 27172
rect 9640 27228 9704 27232
rect 9640 27172 9644 27228
rect 9644 27172 9700 27228
rect 9700 27172 9704 27228
rect 9640 27168 9704 27172
rect 17848 27228 17912 27232
rect 17848 27172 17852 27228
rect 17852 27172 17908 27228
rect 17908 27172 17912 27228
rect 17848 27168 17912 27172
rect 17928 27228 17992 27232
rect 17928 27172 17932 27228
rect 17932 27172 17988 27228
rect 17988 27172 17992 27228
rect 17928 27168 17992 27172
rect 18008 27228 18072 27232
rect 18008 27172 18012 27228
rect 18012 27172 18068 27228
rect 18068 27172 18072 27228
rect 18008 27168 18072 27172
rect 18088 27228 18152 27232
rect 18088 27172 18092 27228
rect 18092 27172 18148 27228
rect 18148 27172 18152 27228
rect 18088 27168 18152 27172
rect 26296 27228 26360 27232
rect 26296 27172 26300 27228
rect 26300 27172 26356 27228
rect 26356 27172 26360 27228
rect 26296 27168 26360 27172
rect 26376 27228 26440 27232
rect 26376 27172 26380 27228
rect 26380 27172 26436 27228
rect 26436 27172 26440 27228
rect 26376 27168 26440 27172
rect 26456 27228 26520 27232
rect 26456 27172 26460 27228
rect 26460 27172 26516 27228
rect 26516 27172 26520 27228
rect 26456 27168 26520 27172
rect 26536 27228 26600 27232
rect 26536 27172 26540 27228
rect 26540 27172 26596 27228
rect 26596 27172 26600 27228
rect 26536 27168 26600 27172
rect 5176 26684 5240 26688
rect 5176 26628 5180 26684
rect 5180 26628 5236 26684
rect 5236 26628 5240 26684
rect 5176 26624 5240 26628
rect 5256 26684 5320 26688
rect 5256 26628 5260 26684
rect 5260 26628 5316 26684
rect 5316 26628 5320 26684
rect 5256 26624 5320 26628
rect 5336 26684 5400 26688
rect 5336 26628 5340 26684
rect 5340 26628 5396 26684
rect 5396 26628 5400 26684
rect 5336 26624 5400 26628
rect 5416 26684 5480 26688
rect 5416 26628 5420 26684
rect 5420 26628 5476 26684
rect 5476 26628 5480 26684
rect 5416 26624 5480 26628
rect 13624 26684 13688 26688
rect 13624 26628 13628 26684
rect 13628 26628 13684 26684
rect 13684 26628 13688 26684
rect 13624 26624 13688 26628
rect 13704 26684 13768 26688
rect 13704 26628 13708 26684
rect 13708 26628 13764 26684
rect 13764 26628 13768 26684
rect 13704 26624 13768 26628
rect 13784 26684 13848 26688
rect 13784 26628 13788 26684
rect 13788 26628 13844 26684
rect 13844 26628 13848 26684
rect 13784 26624 13848 26628
rect 13864 26684 13928 26688
rect 13864 26628 13868 26684
rect 13868 26628 13924 26684
rect 13924 26628 13928 26684
rect 13864 26624 13928 26628
rect 22072 26684 22136 26688
rect 22072 26628 22076 26684
rect 22076 26628 22132 26684
rect 22132 26628 22136 26684
rect 22072 26624 22136 26628
rect 22152 26684 22216 26688
rect 22152 26628 22156 26684
rect 22156 26628 22212 26684
rect 22212 26628 22216 26684
rect 22152 26624 22216 26628
rect 22232 26684 22296 26688
rect 22232 26628 22236 26684
rect 22236 26628 22292 26684
rect 22292 26628 22296 26684
rect 22232 26624 22296 26628
rect 22312 26684 22376 26688
rect 22312 26628 22316 26684
rect 22316 26628 22372 26684
rect 22372 26628 22376 26684
rect 22312 26624 22376 26628
rect 30520 26684 30584 26688
rect 30520 26628 30524 26684
rect 30524 26628 30580 26684
rect 30580 26628 30584 26684
rect 30520 26624 30584 26628
rect 30600 26684 30664 26688
rect 30600 26628 30604 26684
rect 30604 26628 30660 26684
rect 30660 26628 30664 26684
rect 30600 26624 30664 26628
rect 30680 26684 30744 26688
rect 30680 26628 30684 26684
rect 30684 26628 30740 26684
rect 30740 26628 30744 26684
rect 30680 26624 30744 26628
rect 30760 26684 30824 26688
rect 30760 26628 30764 26684
rect 30764 26628 30820 26684
rect 30820 26628 30824 26684
rect 30760 26624 30824 26628
rect 9400 26140 9464 26144
rect 9400 26084 9404 26140
rect 9404 26084 9460 26140
rect 9460 26084 9464 26140
rect 9400 26080 9464 26084
rect 9480 26140 9544 26144
rect 9480 26084 9484 26140
rect 9484 26084 9540 26140
rect 9540 26084 9544 26140
rect 9480 26080 9544 26084
rect 9560 26140 9624 26144
rect 9560 26084 9564 26140
rect 9564 26084 9620 26140
rect 9620 26084 9624 26140
rect 9560 26080 9624 26084
rect 9640 26140 9704 26144
rect 9640 26084 9644 26140
rect 9644 26084 9700 26140
rect 9700 26084 9704 26140
rect 9640 26080 9704 26084
rect 17848 26140 17912 26144
rect 17848 26084 17852 26140
rect 17852 26084 17908 26140
rect 17908 26084 17912 26140
rect 17848 26080 17912 26084
rect 17928 26140 17992 26144
rect 17928 26084 17932 26140
rect 17932 26084 17988 26140
rect 17988 26084 17992 26140
rect 17928 26080 17992 26084
rect 18008 26140 18072 26144
rect 18008 26084 18012 26140
rect 18012 26084 18068 26140
rect 18068 26084 18072 26140
rect 18008 26080 18072 26084
rect 18088 26140 18152 26144
rect 18088 26084 18092 26140
rect 18092 26084 18148 26140
rect 18148 26084 18152 26140
rect 18088 26080 18152 26084
rect 26296 26140 26360 26144
rect 26296 26084 26300 26140
rect 26300 26084 26356 26140
rect 26356 26084 26360 26140
rect 26296 26080 26360 26084
rect 26376 26140 26440 26144
rect 26376 26084 26380 26140
rect 26380 26084 26436 26140
rect 26436 26084 26440 26140
rect 26376 26080 26440 26084
rect 26456 26140 26520 26144
rect 26456 26084 26460 26140
rect 26460 26084 26516 26140
rect 26516 26084 26520 26140
rect 26456 26080 26520 26084
rect 26536 26140 26600 26144
rect 26536 26084 26540 26140
rect 26540 26084 26596 26140
rect 26596 26084 26600 26140
rect 26536 26080 26600 26084
rect 5176 25596 5240 25600
rect 5176 25540 5180 25596
rect 5180 25540 5236 25596
rect 5236 25540 5240 25596
rect 5176 25536 5240 25540
rect 5256 25596 5320 25600
rect 5256 25540 5260 25596
rect 5260 25540 5316 25596
rect 5316 25540 5320 25596
rect 5256 25536 5320 25540
rect 5336 25596 5400 25600
rect 5336 25540 5340 25596
rect 5340 25540 5396 25596
rect 5396 25540 5400 25596
rect 5336 25536 5400 25540
rect 5416 25596 5480 25600
rect 5416 25540 5420 25596
rect 5420 25540 5476 25596
rect 5476 25540 5480 25596
rect 5416 25536 5480 25540
rect 13624 25596 13688 25600
rect 13624 25540 13628 25596
rect 13628 25540 13684 25596
rect 13684 25540 13688 25596
rect 13624 25536 13688 25540
rect 13704 25596 13768 25600
rect 13704 25540 13708 25596
rect 13708 25540 13764 25596
rect 13764 25540 13768 25596
rect 13704 25536 13768 25540
rect 13784 25596 13848 25600
rect 13784 25540 13788 25596
rect 13788 25540 13844 25596
rect 13844 25540 13848 25596
rect 13784 25536 13848 25540
rect 13864 25596 13928 25600
rect 13864 25540 13868 25596
rect 13868 25540 13924 25596
rect 13924 25540 13928 25596
rect 13864 25536 13928 25540
rect 22072 25596 22136 25600
rect 22072 25540 22076 25596
rect 22076 25540 22132 25596
rect 22132 25540 22136 25596
rect 22072 25536 22136 25540
rect 22152 25596 22216 25600
rect 22152 25540 22156 25596
rect 22156 25540 22212 25596
rect 22212 25540 22216 25596
rect 22152 25536 22216 25540
rect 22232 25596 22296 25600
rect 22232 25540 22236 25596
rect 22236 25540 22292 25596
rect 22292 25540 22296 25596
rect 22232 25536 22296 25540
rect 22312 25596 22376 25600
rect 22312 25540 22316 25596
rect 22316 25540 22372 25596
rect 22372 25540 22376 25596
rect 22312 25536 22376 25540
rect 30520 25596 30584 25600
rect 30520 25540 30524 25596
rect 30524 25540 30580 25596
rect 30580 25540 30584 25596
rect 30520 25536 30584 25540
rect 30600 25596 30664 25600
rect 30600 25540 30604 25596
rect 30604 25540 30660 25596
rect 30660 25540 30664 25596
rect 30600 25536 30664 25540
rect 30680 25596 30744 25600
rect 30680 25540 30684 25596
rect 30684 25540 30740 25596
rect 30740 25540 30744 25596
rect 30680 25536 30744 25540
rect 30760 25596 30824 25600
rect 30760 25540 30764 25596
rect 30764 25540 30820 25596
rect 30820 25540 30824 25596
rect 30760 25536 30824 25540
rect 9400 25052 9464 25056
rect 9400 24996 9404 25052
rect 9404 24996 9460 25052
rect 9460 24996 9464 25052
rect 9400 24992 9464 24996
rect 9480 25052 9544 25056
rect 9480 24996 9484 25052
rect 9484 24996 9540 25052
rect 9540 24996 9544 25052
rect 9480 24992 9544 24996
rect 9560 25052 9624 25056
rect 9560 24996 9564 25052
rect 9564 24996 9620 25052
rect 9620 24996 9624 25052
rect 9560 24992 9624 24996
rect 9640 25052 9704 25056
rect 9640 24996 9644 25052
rect 9644 24996 9700 25052
rect 9700 24996 9704 25052
rect 9640 24992 9704 24996
rect 17848 25052 17912 25056
rect 17848 24996 17852 25052
rect 17852 24996 17908 25052
rect 17908 24996 17912 25052
rect 17848 24992 17912 24996
rect 17928 25052 17992 25056
rect 17928 24996 17932 25052
rect 17932 24996 17988 25052
rect 17988 24996 17992 25052
rect 17928 24992 17992 24996
rect 18008 25052 18072 25056
rect 18008 24996 18012 25052
rect 18012 24996 18068 25052
rect 18068 24996 18072 25052
rect 18008 24992 18072 24996
rect 18088 25052 18152 25056
rect 18088 24996 18092 25052
rect 18092 24996 18148 25052
rect 18148 24996 18152 25052
rect 18088 24992 18152 24996
rect 26296 25052 26360 25056
rect 26296 24996 26300 25052
rect 26300 24996 26356 25052
rect 26356 24996 26360 25052
rect 26296 24992 26360 24996
rect 26376 25052 26440 25056
rect 26376 24996 26380 25052
rect 26380 24996 26436 25052
rect 26436 24996 26440 25052
rect 26376 24992 26440 24996
rect 26456 25052 26520 25056
rect 26456 24996 26460 25052
rect 26460 24996 26516 25052
rect 26516 24996 26520 25052
rect 26456 24992 26520 24996
rect 26536 25052 26600 25056
rect 26536 24996 26540 25052
rect 26540 24996 26596 25052
rect 26596 24996 26600 25052
rect 26536 24992 26600 24996
rect 5176 24508 5240 24512
rect 5176 24452 5180 24508
rect 5180 24452 5236 24508
rect 5236 24452 5240 24508
rect 5176 24448 5240 24452
rect 5256 24508 5320 24512
rect 5256 24452 5260 24508
rect 5260 24452 5316 24508
rect 5316 24452 5320 24508
rect 5256 24448 5320 24452
rect 5336 24508 5400 24512
rect 5336 24452 5340 24508
rect 5340 24452 5396 24508
rect 5396 24452 5400 24508
rect 5336 24448 5400 24452
rect 5416 24508 5480 24512
rect 5416 24452 5420 24508
rect 5420 24452 5476 24508
rect 5476 24452 5480 24508
rect 5416 24448 5480 24452
rect 13624 24508 13688 24512
rect 13624 24452 13628 24508
rect 13628 24452 13684 24508
rect 13684 24452 13688 24508
rect 13624 24448 13688 24452
rect 13704 24508 13768 24512
rect 13704 24452 13708 24508
rect 13708 24452 13764 24508
rect 13764 24452 13768 24508
rect 13704 24448 13768 24452
rect 13784 24508 13848 24512
rect 13784 24452 13788 24508
rect 13788 24452 13844 24508
rect 13844 24452 13848 24508
rect 13784 24448 13848 24452
rect 13864 24508 13928 24512
rect 13864 24452 13868 24508
rect 13868 24452 13924 24508
rect 13924 24452 13928 24508
rect 13864 24448 13928 24452
rect 22072 24508 22136 24512
rect 22072 24452 22076 24508
rect 22076 24452 22132 24508
rect 22132 24452 22136 24508
rect 22072 24448 22136 24452
rect 22152 24508 22216 24512
rect 22152 24452 22156 24508
rect 22156 24452 22212 24508
rect 22212 24452 22216 24508
rect 22152 24448 22216 24452
rect 22232 24508 22296 24512
rect 22232 24452 22236 24508
rect 22236 24452 22292 24508
rect 22292 24452 22296 24508
rect 22232 24448 22296 24452
rect 22312 24508 22376 24512
rect 22312 24452 22316 24508
rect 22316 24452 22372 24508
rect 22372 24452 22376 24508
rect 22312 24448 22376 24452
rect 30520 24508 30584 24512
rect 30520 24452 30524 24508
rect 30524 24452 30580 24508
rect 30580 24452 30584 24508
rect 30520 24448 30584 24452
rect 30600 24508 30664 24512
rect 30600 24452 30604 24508
rect 30604 24452 30660 24508
rect 30660 24452 30664 24508
rect 30600 24448 30664 24452
rect 30680 24508 30744 24512
rect 30680 24452 30684 24508
rect 30684 24452 30740 24508
rect 30740 24452 30744 24508
rect 30680 24448 30744 24452
rect 30760 24508 30824 24512
rect 30760 24452 30764 24508
rect 30764 24452 30820 24508
rect 30820 24452 30824 24508
rect 30760 24448 30824 24452
rect 9400 23964 9464 23968
rect 9400 23908 9404 23964
rect 9404 23908 9460 23964
rect 9460 23908 9464 23964
rect 9400 23904 9464 23908
rect 9480 23964 9544 23968
rect 9480 23908 9484 23964
rect 9484 23908 9540 23964
rect 9540 23908 9544 23964
rect 9480 23904 9544 23908
rect 9560 23964 9624 23968
rect 9560 23908 9564 23964
rect 9564 23908 9620 23964
rect 9620 23908 9624 23964
rect 9560 23904 9624 23908
rect 9640 23964 9704 23968
rect 9640 23908 9644 23964
rect 9644 23908 9700 23964
rect 9700 23908 9704 23964
rect 9640 23904 9704 23908
rect 17848 23964 17912 23968
rect 17848 23908 17852 23964
rect 17852 23908 17908 23964
rect 17908 23908 17912 23964
rect 17848 23904 17912 23908
rect 17928 23964 17992 23968
rect 17928 23908 17932 23964
rect 17932 23908 17988 23964
rect 17988 23908 17992 23964
rect 17928 23904 17992 23908
rect 18008 23964 18072 23968
rect 18008 23908 18012 23964
rect 18012 23908 18068 23964
rect 18068 23908 18072 23964
rect 18008 23904 18072 23908
rect 18088 23964 18152 23968
rect 18088 23908 18092 23964
rect 18092 23908 18148 23964
rect 18148 23908 18152 23964
rect 18088 23904 18152 23908
rect 26296 23964 26360 23968
rect 26296 23908 26300 23964
rect 26300 23908 26356 23964
rect 26356 23908 26360 23964
rect 26296 23904 26360 23908
rect 26376 23964 26440 23968
rect 26376 23908 26380 23964
rect 26380 23908 26436 23964
rect 26436 23908 26440 23964
rect 26376 23904 26440 23908
rect 26456 23964 26520 23968
rect 26456 23908 26460 23964
rect 26460 23908 26516 23964
rect 26516 23908 26520 23964
rect 26456 23904 26520 23908
rect 26536 23964 26600 23968
rect 26536 23908 26540 23964
rect 26540 23908 26596 23964
rect 26596 23908 26600 23964
rect 26536 23904 26600 23908
rect 5176 23420 5240 23424
rect 5176 23364 5180 23420
rect 5180 23364 5236 23420
rect 5236 23364 5240 23420
rect 5176 23360 5240 23364
rect 5256 23420 5320 23424
rect 5256 23364 5260 23420
rect 5260 23364 5316 23420
rect 5316 23364 5320 23420
rect 5256 23360 5320 23364
rect 5336 23420 5400 23424
rect 5336 23364 5340 23420
rect 5340 23364 5396 23420
rect 5396 23364 5400 23420
rect 5336 23360 5400 23364
rect 5416 23420 5480 23424
rect 5416 23364 5420 23420
rect 5420 23364 5476 23420
rect 5476 23364 5480 23420
rect 5416 23360 5480 23364
rect 13624 23420 13688 23424
rect 13624 23364 13628 23420
rect 13628 23364 13684 23420
rect 13684 23364 13688 23420
rect 13624 23360 13688 23364
rect 13704 23420 13768 23424
rect 13704 23364 13708 23420
rect 13708 23364 13764 23420
rect 13764 23364 13768 23420
rect 13704 23360 13768 23364
rect 13784 23420 13848 23424
rect 13784 23364 13788 23420
rect 13788 23364 13844 23420
rect 13844 23364 13848 23420
rect 13784 23360 13848 23364
rect 13864 23420 13928 23424
rect 13864 23364 13868 23420
rect 13868 23364 13924 23420
rect 13924 23364 13928 23420
rect 13864 23360 13928 23364
rect 22072 23420 22136 23424
rect 22072 23364 22076 23420
rect 22076 23364 22132 23420
rect 22132 23364 22136 23420
rect 22072 23360 22136 23364
rect 22152 23420 22216 23424
rect 22152 23364 22156 23420
rect 22156 23364 22212 23420
rect 22212 23364 22216 23420
rect 22152 23360 22216 23364
rect 22232 23420 22296 23424
rect 22232 23364 22236 23420
rect 22236 23364 22292 23420
rect 22292 23364 22296 23420
rect 22232 23360 22296 23364
rect 22312 23420 22376 23424
rect 22312 23364 22316 23420
rect 22316 23364 22372 23420
rect 22372 23364 22376 23420
rect 22312 23360 22376 23364
rect 30520 23420 30584 23424
rect 30520 23364 30524 23420
rect 30524 23364 30580 23420
rect 30580 23364 30584 23420
rect 30520 23360 30584 23364
rect 30600 23420 30664 23424
rect 30600 23364 30604 23420
rect 30604 23364 30660 23420
rect 30660 23364 30664 23420
rect 30600 23360 30664 23364
rect 30680 23420 30744 23424
rect 30680 23364 30684 23420
rect 30684 23364 30740 23420
rect 30740 23364 30744 23420
rect 30680 23360 30744 23364
rect 30760 23420 30824 23424
rect 30760 23364 30764 23420
rect 30764 23364 30820 23420
rect 30820 23364 30824 23420
rect 30760 23360 30824 23364
rect 9400 22876 9464 22880
rect 9400 22820 9404 22876
rect 9404 22820 9460 22876
rect 9460 22820 9464 22876
rect 9400 22816 9464 22820
rect 9480 22876 9544 22880
rect 9480 22820 9484 22876
rect 9484 22820 9540 22876
rect 9540 22820 9544 22876
rect 9480 22816 9544 22820
rect 9560 22876 9624 22880
rect 9560 22820 9564 22876
rect 9564 22820 9620 22876
rect 9620 22820 9624 22876
rect 9560 22816 9624 22820
rect 9640 22876 9704 22880
rect 9640 22820 9644 22876
rect 9644 22820 9700 22876
rect 9700 22820 9704 22876
rect 9640 22816 9704 22820
rect 17848 22876 17912 22880
rect 17848 22820 17852 22876
rect 17852 22820 17908 22876
rect 17908 22820 17912 22876
rect 17848 22816 17912 22820
rect 17928 22876 17992 22880
rect 17928 22820 17932 22876
rect 17932 22820 17988 22876
rect 17988 22820 17992 22876
rect 17928 22816 17992 22820
rect 18008 22876 18072 22880
rect 18008 22820 18012 22876
rect 18012 22820 18068 22876
rect 18068 22820 18072 22876
rect 18008 22816 18072 22820
rect 18088 22876 18152 22880
rect 18088 22820 18092 22876
rect 18092 22820 18148 22876
rect 18148 22820 18152 22876
rect 18088 22816 18152 22820
rect 26296 22876 26360 22880
rect 26296 22820 26300 22876
rect 26300 22820 26356 22876
rect 26356 22820 26360 22876
rect 26296 22816 26360 22820
rect 26376 22876 26440 22880
rect 26376 22820 26380 22876
rect 26380 22820 26436 22876
rect 26436 22820 26440 22876
rect 26376 22816 26440 22820
rect 26456 22876 26520 22880
rect 26456 22820 26460 22876
rect 26460 22820 26516 22876
rect 26516 22820 26520 22876
rect 26456 22816 26520 22820
rect 26536 22876 26600 22880
rect 26536 22820 26540 22876
rect 26540 22820 26596 22876
rect 26596 22820 26600 22876
rect 26536 22816 26600 22820
rect 5176 22332 5240 22336
rect 5176 22276 5180 22332
rect 5180 22276 5236 22332
rect 5236 22276 5240 22332
rect 5176 22272 5240 22276
rect 5256 22332 5320 22336
rect 5256 22276 5260 22332
rect 5260 22276 5316 22332
rect 5316 22276 5320 22332
rect 5256 22272 5320 22276
rect 5336 22332 5400 22336
rect 5336 22276 5340 22332
rect 5340 22276 5396 22332
rect 5396 22276 5400 22332
rect 5336 22272 5400 22276
rect 5416 22332 5480 22336
rect 5416 22276 5420 22332
rect 5420 22276 5476 22332
rect 5476 22276 5480 22332
rect 5416 22272 5480 22276
rect 13624 22332 13688 22336
rect 13624 22276 13628 22332
rect 13628 22276 13684 22332
rect 13684 22276 13688 22332
rect 13624 22272 13688 22276
rect 13704 22332 13768 22336
rect 13704 22276 13708 22332
rect 13708 22276 13764 22332
rect 13764 22276 13768 22332
rect 13704 22272 13768 22276
rect 13784 22332 13848 22336
rect 13784 22276 13788 22332
rect 13788 22276 13844 22332
rect 13844 22276 13848 22332
rect 13784 22272 13848 22276
rect 13864 22332 13928 22336
rect 13864 22276 13868 22332
rect 13868 22276 13924 22332
rect 13924 22276 13928 22332
rect 13864 22272 13928 22276
rect 22072 22332 22136 22336
rect 22072 22276 22076 22332
rect 22076 22276 22132 22332
rect 22132 22276 22136 22332
rect 22072 22272 22136 22276
rect 22152 22332 22216 22336
rect 22152 22276 22156 22332
rect 22156 22276 22212 22332
rect 22212 22276 22216 22332
rect 22152 22272 22216 22276
rect 22232 22332 22296 22336
rect 22232 22276 22236 22332
rect 22236 22276 22292 22332
rect 22292 22276 22296 22332
rect 22232 22272 22296 22276
rect 22312 22332 22376 22336
rect 22312 22276 22316 22332
rect 22316 22276 22372 22332
rect 22372 22276 22376 22332
rect 22312 22272 22376 22276
rect 30520 22332 30584 22336
rect 30520 22276 30524 22332
rect 30524 22276 30580 22332
rect 30580 22276 30584 22332
rect 30520 22272 30584 22276
rect 30600 22332 30664 22336
rect 30600 22276 30604 22332
rect 30604 22276 30660 22332
rect 30660 22276 30664 22332
rect 30600 22272 30664 22276
rect 30680 22332 30744 22336
rect 30680 22276 30684 22332
rect 30684 22276 30740 22332
rect 30740 22276 30744 22332
rect 30680 22272 30744 22276
rect 30760 22332 30824 22336
rect 30760 22276 30764 22332
rect 30764 22276 30820 22332
rect 30820 22276 30824 22332
rect 30760 22272 30824 22276
rect 9400 21788 9464 21792
rect 9400 21732 9404 21788
rect 9404 21732 9460 21788
rect 9460 21732 9464 21788
rect 9400 21728 9464 21732
rect 9480 21788 9544 21792
rect 9480 21732 9484 21788
rect 9484 21732 9540 21788
rect 9540 21732 9544 21788
rect 9480 21728 9544 21732
rect 9560 21788 9624 21792
rect 9560 21732 9564 21788
rect 9564 21732 9620 21788
rect 9620 21732 9624 21788
rect 9560 21728 9624 21732
rect 9640 21788 9704 21792
rect 9640 21732 9644 21788
rect 9644 21732 9700 21788
rect 9700 21732 9704 21788
rect 9640 21728 9704 21732
rect 17848 21788 17912 21792
rect 17848 21732 17852 21788
rect 17852 21732 17908 21788
rect 17908 21732 17912 21788
rect 17848 21728 17912 21732
rect 17928 21788 17992 21792
rect 17928 21732 17932 21788
rect 17932 21732 17988 21788
rect 17988 21732 17992 21788
rect 17928 21728 17992 21732
rect 18008 21788 18072 21792
rect 18008 21732 18012 21788
rect 18012 21732 18068 21788
rect 18068 21732 18072 21788
rect 18008 21728 18072 21732
rect 18088 21788 18152 21792
rect 18088 21732 18092 21788
rect 18092 21732 18148 21788
rect 18148 21732 18152 21788
rect 18088 21728 18152 21732
rect 26296 21788 26360 21792
rect 26296 21732 26300 21788
rect 26300 21732 26356 21788
rect 26356 21732 26360 21788
rect 26296 21728 26360 21732
rect 26376 21788 26440 21792
rect 26376 21732 26380 21788
rect 26380 21732 26436 21788
rect 26436 21732 26440 21788
rect 26376 21728 26440 21732
rect 26456 21788 26520 21792
rect 26456 21732 26460 21788
rect 26460 21732 26516 21788
rect 26516 21732 26520 21788
rect 26456 21728 26520 21732
rect 26536 21788 26600 21792
rect 26536 21732 26540 21788
rect 26540 21732 26596 21788
rect 26596 21732 26600 21788
rect 26536 21728 26600 21732
rect 5176 21244 5240 21248
rect 5176 21188 5180 21244
rect 5180 21188 5236 21244
rect 5236 21188 5240 21244
rect 5176 21184 5240 21188
rect 5256 21244 5320 21248
rect 5256 21188 5260 21244
rect 5260 21188 5316 21244
rect 5316 21188 5320 21244
rect 5256 21184 5320 21188
rect 5336 21244 5400 21248
rect 5336 21188 5340 21244
rect 5340 21188 5396 21244
rect 5396 21188 5400 21244
rect 5336 21184 5400 21188
rect 5416 21244 5480 21248
rect 5416 21188 5420 21244
rect 5420 21188 5476 21244
rect 5476 21188 5480 21244
rect 5416 21184 5480 21188
rect 13624 21244 13688 21248
rect 13624 21188 13628 21244
rect 13628 21188 13684 21244
rect 13684 21188 13688 21244
rect 13624 21184 13688 21188
rect 13704 21244 13768 21248
rect 13704 21188 13708 21244
rect 13708 21188 13764 21244
rect 13764 21188 13768 21244
rect 13704 21184 13768 21188
rect 13784 21244 13848 21248
rect 13784 21188 13788 21244
rect 13788 21188 13844 21244
rect 13844 21188 13848 21244
rect 13784 21184 13848 21188
rect 13864 21244 13928 21248
rect 13864 21188 13868 21244
rect 13868 21188 13924 21244
rect 13924 21188 13928 21244
rect 13864 21184 13928 21188
rect 22072 21244 22136 21248
rect 22072 21188 22076 21244
rect 22076 21188 22132 21244
rect 22132 21188 22136 21244
rect 22072 21184 22136 21188
rect 22152 21244 22216 21248
rect 22152 21188 22156 21244
rect 22156 21188 22212 21244
rect 22212 21188 22216 21244
rect 22152 21184 22216 21188
rect 22232 21244 22296 21248
rect 22232 21188 22236 21244
rect 22236 21188 22292 21244
rect 22292 21188 22296 21244
rect 22232 21184 22296 21188
rect 22312 21244 22376 21248
rect 22312 21188 22316 21244
rect 22316 21188 22372 21244
rect 22372 21188 22376 21244
rect 22312 21184 22376 21188
rect 30520 21244 30584 21248
rect 30520 21188 30524 21244
rect 30524 21188 30580 21244
rect 30580 21188 30584 21244
rect 30520 21184 30584 21188
rect 30600 21244 30664 21248
rect 30600 21188 30604 21244
rect 30604 21188 30660 21244
rect 30660 21188 30664 21244
rect 30600 21184 30664 21188
rect 30680 21244 30744 21248
rect 30680 21188 30684 21244
rect 30684 21188 30740 21244
rect 30740 21188 30744 21244
rect 30680 21184 30744 21188
rect 30760 21244 30824 21248
rect 30760 21188 30764 21244
rect 30764 21188 30820 21244
rect 30820 21188 30824 21244
rect 30760 21184 30824 21188
rect 9400 20700 9464 20704
rect 9400 20644 9404 20700
rect 9404 20644 9460 20700
rect 9460 20644 9464 20700
rect 9400 20640 9464 20644
rect 9480 20700 9544 20704
rect 9480 20644 9484 20700
rect 9484 20644 9540 20700
rect 9540 20644 9544 20700
rect 9480 20640 9544 20644
rect 9560 20700 9624 20704
rect 9560 20644 9564 20700
rect 9564 20644 9620 20700
rect 9620 20644 9624 20700
rect 9560 20640 9624 20644
rect 9640 20700 9704 20704
rect 9640 20644 9644 20700
rect 9644 20644 9700 20700
rect 9700 20644 9704 20700
rect 9640 20640 9704 20644
rect 17848 20700 17912 20704
rect 17848 20644 17852 20700
rect 17852 20644 17908 20700
rect 17908 20644 17912 20700
rect 17848 20640 17912 20644
rect 17928 20700 17992 20704
rect 17928 20644 17932 20700
rect 17932 20644 17988 20700
rect 17988 20644 17992 20700
rect 17928 20640 17992 20644
rect 18008 20700 18072 20704
rect 18008 20644 18012 20700
rect 18012 20644 18068 20700
rect 18068 20644 18072 20700
rect 18008 20640 18072 20644
rect 18088 20700 18152 20704
rect 18088 20644 18092 20700
rect 18092 20644 18148 20700
rect 18148 20644 18152 20700
rect 18088 20640 18152 20644
rect 26296 20700 26360 20704
rect 26296 20644 26300 20700
rect 26300 20644 26356 20700
rect 26356 20644 26360 20700
rect 26296 20640 26360 20644
rect 26376 20700 26440 20704
rect 26376 20644 26380 20700
rect 26380 20644 26436 20700
rect 26436 20644 26440 20700
rect 26376 20640 26440 20644
rect 26456 20700 26520 20704
rect 26456 20644 26460 20700
rect 26460 20644 26516 20700
rect 26516 20644 26520 20700
rect 26456 20640 26520 20644
rect 26536 20700 26600 20704
rect 26536 20644 26540 20700
rect 26540 20644 26596 20700
rect 26596 20644 26600 20700
rect 26536 20640 26600 20644
rect 5176 20156 5240 20160
rect 5176 20100 5180 20156
rect 5180 20100 5236 20156
rect 5236 20100 5240 20156
rect 5176 20096 5240 20100
rect 5256 20156 5320 20160
rect 5256 20100 5260 20156
rect 5260 20100 5316 20156
rect 5316 20100 5320 20156
rect 5256 20096 5320 20100
rect 5336 20156 5400 20160
rect 5336 20100 5340 20156
rect 5340 20100 5396 20156
rect 5396 20100 5400 20156
rect 5336 20096 5400 20100
rect 5416 20156 5480 20160
rect 5416 20100 5420 20156
rect 5420 20100 5476 20156
rect 5476 20100 5480 20156
rect 5416 20096 5480 20100
rect 13624 20156 13688 20160
rect 13624 20100 13628 20156
rect 13628 20100 13684 20156
rect 13684 20100 13688 20156
rect 13624 20096 13688 20100
rect 13704 20156 13768 20160
rect 13704 20100 13708 20156
rect 13708 20100 13764 20156
rect 13764 20100 13768 20156
rect 13704 20096 13768 20100
rect 13784 20156 13848 20160
rect 13784 20100 13788 20156
rect 13788 20100 13844 20156
rect 13844 20100 13848 20156
rect 13784 20096 13848 20100
rect 13864 20156 13928 20160
rect 13864 20100 13868 20156
rect 13868 20100 13924 20156
rect 13924 20100 13928 20156
rect 13864 20096 13928 20100
rect 22072 20156 22136 20160
rect 22072 20100 22076 20156
rect 22076 20100 22132 20156
rect 22132 20100 22136 20156
rect 22072 20096 22136 20100
rect 22152 20156 22216 20160
rect 22152 20100 22156 20156
rect 22156 20100 22212 20156
rect 22212 20100 22216 20156
rect 22152 20096 22216 20100
rect 22232 20156 22296 20160
rect 22232 20100 22236 20156
rect 22236 20100 22292 20156
rect 22292 20100 22296 20156
rect 22232 20096 22296 20100
rect 22312 20156 22376 20160
rect 22312 20100 22316 20156
rect 22316 20100 22372 20156
rect 22372 20100 22376 20156
rect 22312 20096 22376 20100
rect 30520 20156 30584 20160
rect 30520 20100 30524 20156
rect 30524 20100 30580 20156
rect 30580 20100 30584 20156
rect 30520 20096 30584 20100
rect 30600 20156 30664 20160
rect 30600 20100 30604 20156
rect 30604 20100 30660 20156
rect 30660 20100 30664 20156
rect 30600 20096 30664 20100
rect 30680 20156 30744 20160
rect 30680 20100 30684 20156
rect 30684 20100 30740 20156
rect 30740 20100 30744 20156
rect 30680 20096 30744 20100
rect 30760 20156 30824 20160
rect 30760 20100 30764 20156
rect 30764 20100 30820 20156
rect 30820 20100 30824 20156
rect 30760 20096 30824 20100
rect 9400 19612 9464 19616
rect 9400 19556 9404 19612
rect 9404 19556 9460 19612
rect 9460 19556 9464 19612
rect 9400 19552 9464 19556
rect 9480 19612 9544 19616
rect 9480 19556 9484 19612
rect 9484 19556 9540 19612
rect 9540 19556 9544 19612
rect 9480 19552 9544 19556
rect 9560 19612 9624 19616
rect 9560 19556 9564 19612
rect 9564 19556 9620 19612
rect 9620 19556 9624 19612
rect 9560 19552 9624 19556
rect 9640 19612 9704 19616
rect 9640 19556 9644 19612
rect 9644 19556 9700 19612
rect 9700 19556 9704 19612
rect 9640 19552 9704 19556
rect 17848 19612 17912 19616
rect 17848 19556 17852 19612
rect 17852 19556 17908 19612
rect 17908 19556 17912 19612
rect 17848 19552 17912 19556
rect 17928 19612 17992 19616
rect 17928 19556 17932 19612
rect 17932 19556 17988 19612
rect 17988 19556 17992 19612
rect 17928 19552 17992 19556
rect 18008 19612 18072 19616
rect 18008 19556 18012 19612
rect 18012 19556 18068 19612
rect 18068 19556 18072 19612
rect 18008 19552 18072 19556
rect 18088 19612 18152 19616
rect 18088 19556 18092 19612
rect 18092 19556 18148 19612
rect 18148 19556 18152 19612
rect 18088 19552 18152 19556
rect 26296 19612 26360 19616
rect 26296 19556 26300 19612
rect 26300 19556 26356 19612
rect 26356 19556 26360 19612
rect 26296 19552 26360 19556
rect 26376 19612 26440 19616
rect 26376 19556 26380 19612
rect 26380 19556 26436 19612
rect 26436 19556 26440 19612
rect 26376 19552 26440 19556
rect 26456 19612 26520 19616
rect 26456 19556 26460 19612
rect 26460 19556 26516 19612
rect 26516 19556 26520 19612
rect 26456 19552 26520 19556
rect 26536 19612 26600 19616
rect 26536 19556 26540 19612
rect 26540 19556 26596 19612
rect 26596 19556 26600 19612
rect 26536 19552 26600 19556
rect 5176 19068 5240 19072
rect 5176 19012 5180 19068
rect 5180 19012 5236 19068
rect 5236 19012 5240 19068
rect 5176 19008 5240 19012
rect 5256 19068 5320 19072
rect 5256 19012 5260 19068
rect 5260 19012 5316 19068
rect 5316 19012 5320 19068
rect 5256 19008 5320 19012
rect 5336 19068 5400 19072
rect 5336 19012 5340 19068
rect 5340 19012 5396 19068
rect 5396 19012 5400 19068
rect 5336 19008 5400 19012
rect 5416 19068 5480 19072
rect 5416 19012 5420 19068
rect 5420 19012 5476 19068
rect 5476 19012 5480 19068
rect 5416 19008 5480 19012
rect 13624 19068 13688 19072
rect 13624 19012 13628 19068
rect 13628 19012 13684 19068
rect 13684 19012 13688 19068
rect 13624 19008 13688 19012
rect 13704 19068 13768 19072
rect 13704 19012 13708 19068
rect 13708 19012 13764 19068
rect 13764 19012 13768 19068
rect 13704 19008 13768 19012
rect 13784 19068 13848 19072
rect 13784 19012 13788 19068
rect 13788 19012 13844 19068
rect 13844 19012 13848 19068
rect 13784 19008 13848 19012
rect 13864 19068 13928 19072
rect 13864 19012 13868 19068
rect 13868 19012 13924 19068
rect 13924 19012 13928 19068
rect 13864 19008 13928 19012
rect 22072 19068 22136 19072
rect 22072 19012 22076 19068
rect 22076 19012 22132 19068
rect 22132 19012 22136 19068
rect 22072 19008 22136 19012
rect 22152 19068 22216 19072
rect 22152 19012 22156 19068
rect 22156 19012 22212 19068
rect 22212 19012 22216 19068
rect 22152 19008 22216 19012
rect 22232 19068 22296 19072
rect 22232 19012 22236 19068
rect 22236 19012 22292 19068
rect 22292 19012 22296 19068
rect 22232 19008 22296 19012
rect 22312 19068 22376 19072
rect 22312 19012 22316 19068
rect 22316 19012 22372 19068
rect 22372 19012 22376 19068
rect 22312 19008 22376 19012
rect 30520 19068 30584 19072
rect 30520 19012 30524 19068
rect 30524 19012 30580 19068
rect 30580 19012 30584 19068
rect 30520 19008 30584 19012
rect 30600 19068 30664 19072
rect 30600 19012 30604 19068
rect 30604 19012 30660 19068
rect 30660 19012 30664 19068
rect 30600 19008 30664 19012
rect 30680 19068 30744 19072
rect 30680 19012 30684 19068
rect 30684 19012 30740 19068
rect 30740 19012 30744 19068
rect 30680 19008 30744 19012
rect 30760 19068 30824 19072
rect 30760 19012 30764 19068
rect 30764 19012 30820 19068
rect 30820 19012 30824 19068
rect 30760 19008 30824 19012
rect 9400 18524 9464 18528
rect 9400 18468 9404 18524
rect 9404 18468 9460 18524
rect 9460 18468 9464 18524
rect 9400 18464 9464 18468
rect 9480 18524 9544 18528
rect 9480 18468 9484 18524
rect 9484 18468 9540 18524
rect 9540 18468 9544 18524
rect 9480 18464 9544 18468
rect 9560 18524 9624 18528
rect 9560 18468 9564 18524
rect 9564 18468 9620 18524
rect 9620 18468 9624 18524
rect 9560 18464 9624 18468
rect 9640 18524 9704 18528
rect 9640 18468 9644 18524
rect 9644 18468 9700 18524
rect 9700 18468 9704 18524
rect 9640 18464 9704 18468
rect 17848 18524 17912 18528
rect 17848 18468 17852 18524
rect 17852 18468 17908 18524
rect 17908 18468 17912 18524
rect 17848 18464 17912 18468
rect 17928 18524 17992 18528
rect 17928 18468 17932 18524
rect 17932 18468 17988 18524
rect 17988 18468 17992 18524
rect 17928 18464 17992 18468
rect 18008 18524 18072 18528
rect 18008 18468 18012 18524
rect 18012 18468 18068 18524
rect 18068 18468 18072 18524
rect 18008 18464 18072 18468
rect 18088 18524 18152 18528
rect 18088 18468 18092 18524
rect 18092 18468 18148 18524
rect 18148 18468 18152 18524
rect 18088 18464 18152 18468
rect 26296 18524 26360 18528
rect 26296 18468 26300 18524
rect 26300 18468 26356 18524
rect 26356 18468 26360 18524
rect 26296 18464 26360 18468
rect 26376 18524 26440 18528
rect 26376 18468 26380 18524
rect 26380 18468 26436 18524
rect 26436 18468 26440 18524
rect 26376 18464 26440 18468
rect 26456 18524 26520 18528
rect 26456 18468 26460 18524
rect 26460 18468 26516 18524
rect 26516 18468 26520 18524
rect 26456 18464 26520 18468
rect 26536 18524 26600 18528
rect 26536 18468 26540 18524
rect 26540 18468 26596 18524
rect 26596 18468 26600 18524
rect 26536 18464 26600 18468
rect 5176 17980 5240 17984
rect 5176 17924 5180 17980
rect 5180 17924 5236 17980
rect 5236 17924 5240 17980
rect 5176 17920 5240 17924
rect 5256 17980 5320 17984
rect 5256 17924 5260 17980
rect 5260 17924 5316 17980
rect 5316 17924 5320 17980
rect 5256 17920 5320 17924
rect 5336 17980 5400 17984
rect 5336 17924 5340 17980
rect 5340 17924 5396 17980
rect 5396 17924 5400 17980
rect 5336 17920 5400 17924
rect 5416 17980 5480 17984
rect 5416 17924 5420 17980
rect 5420 17924 5476 17980
rect 5476 17924 5480 17980
rect 5416 17920 5480 17924
rect 13624 17980 13688 17984
rect 13624 17924 13628 17980
rect 13628 17924 13684 17980
rect 13684 17924 13688 17980
rect 13624 17920 13688 17924
rect 13704 17980 13768 17984
rect 13704 17924 13708 17980
rect 13708 17924 13764 17980
rect 13764 17924 13768 17980
rect 13704 17920 13768 17924
rect 13784 17980 13848 17984
rect 13784 17924 13788 17980
rect 13788 17924 13844 17980
rect 13844 17924 13848 17980
rect 13784 17920 13848 17924
rect 13864 17980 13928 17984
rect 13864 17924 13868 17980
rect 13868 17924 13924 17980
rect 13924 17924 13928 17980
rect 13864 17920 13928 17924
rect 22072 17980 22136 17984
rect 22072 17924 22076 17980
rect 22076 17924 22132 17980
rect 22132 17924 22136 17980
rect 22072 17920 22136 17924
rect 22152 17980 22216 17984
rect 22152 17924 22156 17980
rect 22156 17924 22212 17980
rect 22212 17924 22216 17980
rect 22152 17920 22216 17924
rect 22232 17980 22296 17984
rect 22232 17924 22236 17980
rect 22236 17924 22292 17980
rect 22292 17924 22296 17980
rect 22232 17920 22296 17924
rect 22312 17980 22376 17984
rect 22312 17924 22316 17980
rect 22316 17924 22372 17980
rect 22372 17924 22376 17980
rect 22312 17920 22376 17924
rect 30520 17980 30584 17984
rect 30520 17924 30524 17980
rect 30524 17924 30580 17980
rect 30580 17924 30584 17980
rect 30520 17920 30584 17924
rect 30600 17980 30664 17984
rect 30600 17924 30604 17980
rect 30604 17924 30660 17980
rect 30660 17924 30664 17980
rect 30600 17920 30664 17924
rect 30680 17980 30744 17984
rect 30680 17924 30684 17980
rect 30684 17924 30740 17980
rect 30740 17924 30744 17980
rect 30680 17920 30744 17924
rect 30760 17980 30824 17984
rect 30760 17924 30764 17980
rect 30764 17924 30820 17980
rect 30820 17924 30824 17980
rect 30760 17920 30824 17924
rect 9400 17436 9464 17440
rect 9400 17380 9404 17436
rect 9404 17380 9460 17436
rect 9460 17380 9464 17436
rect 9400 17376 9464 17380
rect 9480 17436 9544 17440
rect 9480 17380 9484 17436
rect 9484 17380 9540 17436
rect 9540 17380 9544 17436
rect 9480 17376 9544 17380
rect 9560 17436 9624 17440
rect 9560 17380 9564 17436
rect 9564 17380 9620 17436
rect 9620 17380 9624 17436
rect 9560 17376 9624 17380
rect 9640 17436 9704 17440
rect 9640 17380 9644 17436
rect 9644 17380 9700 17436
rect 9700 17380 9704 17436
rect 9640 17376 9704 17380
rect 17848 17436 17912 17440
rect 17848 17380 17852 17436
rect 17852 17380 17908 17436
rect 17908 17380 17912 17436
rect 17848 17376 17912 17380
rect 17928 17436 17992 17440
rect 17928 17380 17932 17436
rect 17932 17380 17988 17436
rect 17988 17380 17992 17436
rect 17928 17376 17992 17380
rect 18008 17436 18072 17440
rect 18008 17380 18012 17436
rect 18012 17380 18068 17436
rect 18068 17380 18072 17436
rect 18008 17376 18072 17380
rect 18088 17436 18152 17440
rect 18088 17380 18092 17436
rect 18092 17380 18148 17436
rect 18148 17380 18152 17436
rect 18088 17376 18152 17380
rect 26296 17436 26360 17440
rect 26296 17380 26300 17436
rect 26300 17380 26356 17436
rect 26356 17380 26360 17436
rect 26296 17376 26360 17380
rect 26376 17436 26440 17440
rect 26376 17380 26380 17436
rect 26380 17380 26436 17436
rect 26436 17380 26440 17436
rect 26376 17376 26440 17380
rect 26456 17436 26520 17440
rect 26456 17380 26460 17436
rect 26460 17380 26516 17436
rect 26516 17380 26520 17436
rect 26456 17376 26520 17380
rect 26536 17436 26600 17440
rect 26536 17380 26540 17436
rect 26540 17380 26596 17436
rect 26596 17380 26600 17436
rect 26536 17376 26600 17380
rect 5176 16892 5240 16896
rect 5176 16836 5180 16892
rect 5180 16836 5236 16892
rect 5236 16836 5240 16892
rect 5176 16832 5240 16836
rect 5256 16892 5320 16896
rect 5256 16836 5260 16892
rect 5260 16836 5316 16892
rect 5316 16836 5320 16892
rect 5256 16832 5320 16836
rect 5336 16892 5400 16896
rect 5336 16836 5340 16892
rect 5340 16836 5396 16892
rect 5396 16836 5400 16892
rect 5336 16832 5400 16836
rect 5416 16892 5480 16896
rect 5416 16836 5420 16892
rect 5420 16836 5476 16892
rect 5476 16836 5480 16892
rect 5416 16832 5480 16836
rect 13624 16892 13688 16896
rect 13624 16836 13628 16892
rect 13628 16836 13684 16892
rect 13684 16836 13688 16892
rect 13624 16832 13688 16836
rect 13704 16892 13768 16896
rect 13704 16836 13708 16892
rect 13708 16836 13764 16892
rect 13764 16836 13768 16892
rect 13704 16832 13768 16836
rect 13784 16892 13848 16896
rect 13784 16836 13788 16892
rect 13788 16836 13844 16892
rect 13844 16836 13848 16892
rect 13784 16832 13848 16836
rect 13864 16892 13928 16896
rect 13864 16836 13868 16892
rect 13868 16836 13924 16892
rect 13924 16836 13928 16892
rect 13864 16832 13928 16836
rect 22072 16892 22136 16896
rect 22072 16836 22076 16892
rect 22076 16836 22132 16892
rect 22132 16836 22136 16892
rect 22072 16832 22136 16836
rect 22152 16892 22216 16896
rect 22152 16836 22156 16892
rect 22156 16836 22212 16892
rect 22212 16836 22216 16892
rect 22152 16832 22216 16836
rect 22232 16892 22296 16896
rect 22232 16836 22236 16892
rect 22236 16836 22292 16892
rect 22292 16836 22296 16892
rect 22232 16832 22296 16836
rect 22312 16892 22376 16896
rect 22312 16836 22316 16892
rect 22316 16836 22372 16892
rect 22372 16836 22376 16892
rect 22312 16832 22376 16836
rect 30520 16892 30584 16896
rect 30520 16836 30524 16892
rect 30524 16836 30580 16892
rect 30580 16836 30584 16892
rect 30520 16832 30584 16836
rect 30600 16892 30664 16896
rect 30600 16836 30604 16892
rect 30604 16836 30660 16892
rect 30660 16836 30664 16892
rect 30600 16832 30664 16836
rect 30680 16892 30744 16896
rect 30680 16836 30684 16892
rect 30684 16836 30740 16892
rect 30740 16836 30744 16892
rect 30680 16832 30744 16836
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 9400 16348 9464 16352
rect 9400 16292 9404 16348
rect 9404 16292 9460 16348
rect 9460 16292 9464 16348
rect 9400 16288 9464 16292
rect 9480 16348 9544 16352
rect 9480 16292 9484 16348
rect 9484 16292 9540 16348
rect 9540 16292 9544 16348
rect 9480 16288 9544 16292
rect 9560 16348 9624 16352
rect 9560 16292 9564 16348
rect 9564 16292 9620 16348
rect 9620 16292 9624 16348
rect 9560 16288 9624 16292
rect 9640 16348 9704 16352
rect 9640 16292 9644 16348
rect 9644 16292 9700 16348
rect 9700 16292 9704 16348
rect 9640 16288 9704 16292
rect 17848 16348 17912 16352
rect 17848 16292 17852 16348
rect 17852 16292 17908 16348
rect 17908 16292 17912 16348
rect 17848 16288 17912 16292
rect 17928 16348 17992 16352
rect 17928 16292 17932 16348
rect 17932 16292 17988 16348
rect 17988 16292 17992 16348
rect 17928 16288 17992 16292
rect 18008 16348 18072 16352
rect 18008 16292 18012 16348
rect 18012 16292 18068 16348
rect 18068 16292 18072 16348
rect 18008 16288 18072 16292
rect 18088 16348 18152 16352
rect 18088 16292 18092 16348
rect 18092 16292 18148 16348
rect 18148 16292 18152 16348
rect 18088 16288 18152 16292
rect 26296 16348 26360 16352
rect 26296 16292 26300 16348
rect 26300 16292 26356 16348
rect 26356 16292 26360 16348
rect 26296 16288 26360 16292
rect 26376 16348 26440 16352
rect 26376 16292 26380 16348
rect 26380 16292 26436 16348
rect 26436 16292 26440 16348
rect 26376 16288 26440 16292
rect 26456 16348 26520 16352
rect 26456 16292 26460 16348
rect 26460 16292 26516 16348
rect 26516 16292 26520 16348
rect 26456 16288 26520 16292
rect 26536 16348 26600 16352
rect 26536 16292 26540 16348
rect 26540 16292 26596 16348
rect 26596 16292 26600 16348
rect 26536 16288 26600 16292
rect 5176 15804 5240 15808
rect 5176 15748 5180 15804
rect 5180 15748 5236 15804
rect 5236 15748 5240 15804
rect 5176 15744 5240 15748
rect 5256 15804 5320 15808
rect 5256 15748 5260 15804
rect 5260 15748 5316 15804
rect 5316 15748 5320 15804
rect 5256 15744 5320 15748
rect 5336 15804 5400 15808
rect 5336 15748 5340 15804
rect 5340 15748 5396 15804
rect 5396 15748 5400 15804
rect 5336 15744 5400 15748
rect 5416 15804 5480 15808
rect 5416 15748 5420 15804
rect 5420 15748 5476 15804
rect 5476 15748 5480 15804
rect 5416 15744 5480 15748
rect 13624 15804 13688 15808
rect 13624 15748 13628 15804
rect 13628 15748 13684 15804
rect 13684 15748 13688 15804
rect 13624 15744 13688 15748
rect 13704 15804 13768 15808
rect 13704 15748 13708 15804
rect 13708 15748 13764 15804
rect 13764 15748 13768 15804
rect 13704 15744 13768 15748
rect 13784 15804 13848 15808
rect 13784 15748 13788 15804
rect 13788 15748 13844 15804
rect 13844 15748 13848 15804
rect 13784 15744 13848 15748
rect 13864 15804 13928 15808
rect 13864 15748 13868 15804
rect 13868 15748 13924 15804
rect 13924 15748 13928 15804
rect 13864 15744 13928 15748
rect 22072 15804 22136 15808
rect 22072 15748 22076 15804
rect 22076 15748 22132 15804
rect 22132 15748 22136 15804
rect 22072 15744 22136 15748
rect 22152 15804 22216 15808
rect 22152 15748 22156 15804
rect 22156 15748 22212 15804
rect 22212 15748 22216 15804
rect 22152 15744 22216 15748
rect 22232 15804 22296 15808
rect 22232 15748 22236 15804
rect 22236 15748 22292 15804
rect 22292 15748 22296 15804
rect 22232 15744 22296 15748
rect 22312 15804 22376 15808
rect 22312 15748 22316 15804
rect 22316 15748 22372 15804
rect 22372 15748 22376 15804
rect 22312 15744 22376 15748
rect 30520 15804 30584 15808
rect 30520 15748 30524 15804
rect 30524 15748 30580 15804
rect 30580 15748 30584 15804
rect 30520 15744 30584 15748
rect 30600 15804 30664 15808
rect 30600 15748 30604 15804
rect 30604 15748 30660 15804
rect 30660 15748 30664 15804
rect 30600 15744 30664 15748
rect 30680 15804 30744 15808
rect 30680 15748 30684 15804
rect 30684 15748 30740 15804
rect 30740 15748 30744 15804
rect 30680 15744 30744 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 9400 15260 9464 15264
rect 9400 15204 9404 15260
rect 9404 15204 9460 15260
rect 9460 15204 9464 15260
rect 9400 15200 9464 15204
rect 9480 15260 9544 15264
rect 9480 15204 9484 15260
rect 9484 15204 9540 15260
rect 9540 15204 9544 15260
rect 9480 15200 9544 15204
rect 9560 15260 9624 15264
rect 9560 15204 9564 15260
rect 9564 15204 9620 15260
rect 9620 15204 9624 15260
rect 9560 15200 9624 15204
rect 9640 15260 9704 15264
rect 9640 15204 9644 15260
rect 9644 15204 9700 15260
rect 9700 15204 9704 15260
rect 9640 15200 9704 15204
rect 17848 15260 17912 15264
rect 17848 15204 17852 15260
rect 17852 15204 17908 15260
rect 17908 15204 17912 15260
rect 17848 15200 17912 15204
rect 17928 15260 17992 15264
rect 17928 15204 17932 15260
rect 17932 15204 17988 15260
rect 17988 15204 17992 15260
rect 17928 15200 17992 15204
rect 18008 15260 18072 15264
rect 18008 15204 18012 15260
rect 18012 15204 18068 15260
rect 18068 15204 18072 15260
rect 18008 15200 18072 15204
rect 18088 15260 18152 15264
rect 18088 15204 18092 15260
rect 18092 15204 18148 15260
rect 18148 15204 18152 15260
rect 18088 15200 18152 15204
rect 26296 15260 26360 15264
rect 26296 15204 26300 15260
rect 26300 15204 26356 15260
rect 26356 15204 26360 15260
rect 26296 15200 26360 15204
rect 26376 15260 26440 15264
rect 26376 15204 26380 15260
rect 26380 15204 26436 15260
rect 26436 15204 26440 15260
rect 26376 15200 26440 15204
rect 26456 15260 26520 15264
rect 26456 15204 26460 15260
rect 26460 15204 26516 15260
rect 26516 15204 26520 15260
rect 26456 15200 26520 15204
rect 26536 15260 26600 15264
rect 26536 15204 26540 15260
rect 26540 15204 26596 15260
rect 26596 15204 26600 15260
rect 26536 15200 26600 15204
rect 5176 14716 5240 14720
rect 5176 14660 5180 14716
rect 5180 14660 5236 14716
rect 5236 14660 5240 14716
rect 5176 14656 5240 14660
rect 5256 14716 5320 14720
rect 5256 14660 5260 14716
rect 5260 14660 5316 14716
rect 5316 14660 5320 14716
rect 5256 14656 5320 14660
rect 5336 14716 5400 14720
rect 5336 14660 5340 14716
rect 5340 14660 5396 14716
rect 5396 14660 5400 14716
rect 5336 14656 5400 14660
rect 5416 14716 5480 14720
rect 5416 14660 5420 14716
rect 5420 14660 5476 14716
rect 5476 14660 5480 14716
rect 5416 14656 5480 14660
rect 13624 14716 13688 14720
rect 13624 14660 13628 14716
rect 13628 14660 13684 14716
rect 13684 14660 13688 14716
rect 13624 14656 13688 14660
rect 13704 14716 13768 14720
rect 13704 14660 13708 14716
rect 13708 14660 13764 14716
rect 13764 14660 13768 14716
rect 13704 14656 13768 14660
rect 13784 14716 13848 14720
rect 13784 14660 13788 14716
rect 13788 14660 13844 14716
rect 13844 14660 13848 14716
rect 13784 14656 13848 14660
rect 13864 14716 13928 14720
rect 13864 14660 13868 14716
rect 13868 14660 13924 14716
rect 13924 14660 13928 14716
rect 13864 14656 13928 14660
rect 22072 14716 22136 14720
rect 22072 14660 22076 14716
rect 22076 14660 22132 14716
rect 22132 14660 22136 14716
rect 22072 14656 22136 14660
rect 22152 14716 22216 14720
rect 22152 14660 22156 14716
rect 22156 14660 22212 14716
rect 22212 14660 22216 14716
rect 22152 14656 22216 14660
rect 22232 14716 22296 14720
rect 22232 14660 22236 14716
rect 22236 14660 22292 14716
rect 22292 14660 22296 14716
rect 22232 14656 22296 14660
rect 22312 14716 22376 14720
rect 22312 14660 22316 14716
rect 22316 14660 22372 14716
rect 22372 14660 22376 14716
rect 22312 14656 22376 14660
rect 30520 14716 30584 14720
rect 30520 14660 30524 14716
rect 30524 14660 30580 14716
rect 30580 14660 30584 14716
rect 30520 14656 30584 14660
rect 30600 14716 30664 14720
rect 30600 14660 30604 14716
rect 30604 14660 30660 14716
rect 30660 14660 30664 14716
rect 30600 14656 30664 14660
rect 30680 14716 30744 14720
rect 30680 14660 30684 14716
rect 30684 14660 30740 14716
rect 30740 14660 30744 14716
rect 30680 14656 30744 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 9400 14172 9464 14176
rect 9400 14116 9404 14172
rect 9404 14116 9460 14172
rect 9460 14116 9464 14172
rect 9400 14112 9464 14116
rect 9480 14172 9544 14176
rect 9480 14116 9484 14172
rect 9484 14116 9540 14172
rect 9540 14116 9544 14172
rect 9480 14112 9544 14116
rect 9560 14172 9624 14176
rect 9560 14116 9564 14172
rect 9564 14116 9620 14172
rect 9620 14116 9624 14172
rect 9560 14112 9624 14116
rect 9640 14172 9704 14176
rect 9640 14116 9644 14172
rect 9644 14116 9700 14172
rect 9700 14116 9704 14172
rect 9640 14112 9704 14116
rect 17848 14172 17912 14176
rect 17848 14116 17852 14172
rect 17852 14116 17908 14172
rect 17908 14116 17912 14172
rect 17848 14112 17912 14116
rect 17928 14172 17992 14176
rect 17928 14116 17932 14172
rect 17932 14116 17988 14172
rect 17988 14116 17992 14172
rect 17928 14112 17992 14116
rect 18008 14172 18072 14176
rect 18008 14116 18012 14172
rect 18012 14116 18068 14172
rect 18068 14116 18072 14172
rect 18008 14112 18072 14116
rect 18088 14172 18152 14176
rect 18088 14116 18092 14172
rect 18092 14116 18148 14172
rect 18148 14116 18152 14172
rect 18088 14112 18152 14116
rect 26296 14172 26360 14176
rect 26296 14116 26300 14172
rect 26300 14116 26356 14172
rect 26356 14116 26360 14172
rect 26296 14112 26360 14116
rect 26376 14172 26440 14176
rect 26376 14116 26380 14172
rect 26380 14116 26436 14172
rect 26436 14116 26440 14172
rect 26376 14112 26440 14116
rect 26456 14172 26520 14176
rect 26456 14116 26460 14172
rect 26460 14116 26516 14172
rect 26516 14116 26520 14172
rect 26456 14112 26520 14116
rect 26536 14172 26600 14176
rect 26536 14116 26540 14172
rect 26540 14116 26596 14172
rect 26596 14116 26600 14172
rect 26536 14112 26600 14116
rect 5176 13628 5240 13632
rect 5176 13572 5180 13628
rect 5180 13572 5236 13628
rect 5236 13572 5240 13628
rect 5176 13568 5240 13572
rect 5256 13628 5320 13632
rect 5256 13572 5260 13628
rect 5260 13572 5316 13628
rect 5316 13572 5320 13628
rect 5256 13568 5320 13572
rect 5336 13628 5400 13632
rect 5336 13572 5340 13628
rect 5340 13572 5396 13628
rect 5396 13572 5400 13628
rect 5336 13568 5400 13572
rect 5416 13628 5480 13632
rect 5416 13572 5420 13628
rect 5420 13572 5476 13628
rect 5476 13572 5480 13628
rect 5416 13568 5480 13572
rect 13624 13628 13688 13632
rect 13624 13572 13628 13628
rect 13628 13572 13684 13628
rect 13684 13572 13688 13628
rect 13624 13568 13688 13572
rect 13704 13628 13768 13632
rect 13704 13572 13708 13628
rect 13708 13572 13764 13628
rect 13764 13572 13768 13628
rect 13704 13568 13768 13572
rect 13784 13628 13848 13632
rect 13784 13572 13788 13628
rect 13788 13572 13844 13628
rect 13844 13572 13848 13628
rect 13784 13568 13848 13572
rect 13864 13628 13928 13632
rect 13864 13572 13868 13628
rect 13868 13572 13924 13628
rect 13924 13572 13928 13628
rect 13864 13568 13928 13572
rect 22072 13628 22136 13632
rect 22072 13572 22076 13628
rect 22076 13572 22132 13628
rect 22132 13572 22136 13628
rect 22072 13568 22136 13572
rect 22152 13628 22216 13632
rect 22152 13572 22156 13628
rect 22156 13572 22212 13628
rect 22212 13572 22216 13628
rect 22152 13568 22216 13572
rect 22232 13628 22296 13632
rect 22232 13572 22236 13628
rect 22236 13572 22292 13628
rect 22292 13572 22296 13628
rect 22232 13568 22296 13572
rect 22312 13628 22376 13632
rect 22312 13572 22316 13628
rect 22316 13572 22372 13628
rect 22372 13572 22376 13628
rect 22312 13568 22376 13572
rect 30520 13628 30584 13632
rect 30520 13572 30524 13628
rect 30524 13572 30580 13628
rect 30580 13572 30584 13628
rect 30520 13568 30584 13572
rect 30600 13628 30664 13632
rect 30600 13572 30604 13628
rect 30604 13572 30660 13628
rect 30660 13572 30664 13628
rect 30600 13568 30664 13572
rect 30680 13628 30744 13632
rect 30680 13572 30684 13628
rect 30684 13572 30740 13628
rect 30740 13572 30744 13628
rect 30680 13568 30744 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 9400 13084 9464 13088
rect 9400 13028 9404 13084
rect 9404 13028 9460 13084
rect 9460 13028 9464 13084
rect 9400 13024 9464 13028
rect 9480 13084 9544 13088
rect 9480 13028 9484 13084
rect 9484 13028 9540 13084
rect 9540 13028 9544 13084
rect 9480 13024 9544 13028
rect 9560 13084 9624 13088
rect 9560 13028 9564 13084
rect 9564 13028 9620 13084
rect 9620 13028 9624 13084
rect 9560 13024 9624 13028
rect 9640 13084 9704 13088
rect 9640 13028 9644 13084
rect 9644 13028 9700 13084
rect 9700 13028 9704 13084
rect 9640 13024 9704 13028
rect 17848 13084 17912 13088
rect 17848 13028 17852 13084
rect 17852 13028 17908 13084
rect 17908 13028 17912 13084
rect 17848 13024 17912 13028
rect 17928 13084 17992 13088
rect 17928 13028 17932 13084
rect 17932 13028 17988 13084
rect 17988 13028 17992 13084
rect 17928 13024 17992 13028
rect 18008 13084 18072 13088
rect 18008 13028 18012 13084
rect 18012 13028 18068 13084
rect 18068 13028 18072 13084
rect 18008 13024 18072 13028
rect 18088 13084 18152 13088
rect 18088 13028 18092 13084
rect 18092 13028 18148 13084
rect 18148 13028 18152 13084
rect 18088 13024 18152 13028
rect 26296 13084 26360 13088
rect 26296 13028 26300 13084
rect 26300 13028 26356 13084
rect 26356 13028 26360 13084
rect 26296 13024 26360 13028
rect 26376 13084 26440 13088
rect 26376 13028 26380 13084
rect 26380 13028 26436 13084
rect 26436 13028 26440 13084
rect 26376 13024 26440 13028
rect 26456 13084 26520 13088
rect 26456 13028 26460 13084
rect 26460 13028 26516 13084
rect 26516 13028 26520 13084
rect 26456 13024 26520 13028
rect 26536 13084 26600 13088
rect 26536 13028 26540 13084
rect 26540 13028 26596 13084
rect 26596 13028 26600 13084
rect 26536 13024 26600 13028
rect 5176 12540 5240 12544
rect 5176 12484 5180 12540
rect 5180 12484 5236 12540
rect 5236 12484 5240 12540
rect 5176 12480 5240 12484
rect 5256 12540 5320 12544
rect 5256 12484 5260 12540
rect 5260 12484 5316 12540
rect 5316 12484 5320 12540
rect 5256 12480 5320 12484
rect 5336 12540 5400 12544
rect 5336 12484 5340 12540
rect 5340 12484 5396 12540
rect 5396 12484 5400 12540
rect 5336 12480 5400 12484
rect 5416 12540 5480 12544
rect 5416 12484 5420 12540
rect 5420 12484 5476 12540
rect 5476 12484 5480 12540
rect 5416 12480 5480 12484
rect 13624 12540 13688 12544
rect 13624 12484 13628 12540
rect 13628 12484 13684 12540
rect 13684 12484 13688 12540
rect 13624 12480 13688 12484
rect 13704 12540 13768 12544
rect 13704 12484 13708 12540
rect 13708 12484 13764 12540
rect 13764 12484 13768 12540
rect 13704 12480 13768 12484
rect 13784 12540 13848 12544
rect 13784 12484 13788 12540
rect 13788 12484 13844 12540
rect 13844 12484 13848 12540
rect 13784 12480 13848 12484
rect 13864 12540 13928 12544
rect 13864 12484 13868 12540
rect 13868 12484 13924 12540
rect 13924 12484 13928 12540
rect 13864 12480 13928 12484
rect 22072 12540 22136 12544
rect 22072 12484 22076 12540
rect 22076 12484 22132 12540
rect 22132 12484 22136 12540
rect 22072 12480 22136 12484
rect 22152 12540 22216 12544
rect 22152 12484 22156 12540
rect 22156 12484 22212 12540
rect 22212 12484 22216 12540
rect 22152 12480 22216 12484
rect 22232 12540 22296 12544
rect 22232 12484 22236 12540
rect 22236 12484 22292 12540
rect 22292 12484 22296 12540
rect 22232 12480 22296 12484
rect 22312 12540 22376 12544
rect 22312 12484 22316 12540
rect 22316 12484 22372 12540
rect 22372 12484 22376 12540
rect 22312 12480 22376 12484
rect 30520 12540 30584 12544
rect 30520 12484 30524 12540
rect 30524 12484 30580 12540
rect 30580 12484 30584 12540
rect 30520 12480 30584 12484
rect 30600 12540 30664 12544
rect 30600 12484 30604 12540
rect 30604 12484 30660 12540
rect 30660 12484 30664 12540
rect 30600 12480 30664 12484
rect 30680 12540 30744 12544
rect 30680 12484 30684 12540
rect 30684 12484 30740 12540
rect 30740 12484 30744 12540
rect 30680 12480 30744 12484
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 9400 11996 9464 12000
rect 9400 11940 9404 11996
rect 9404 11940 9460 11996
rect 9460 11940 9464 11996
rect 9400 11936 9464 11940
rect 9480 11996 9544 12000
rect 9480 11940 9484 11996
rect 9484 11940 9540 11996
rect 9540 11940 9544 11996
rect 9480 11936 9544 11940
rect 9560 11996 9624 12000
rect 9560 11940 9564 11996
rect 9564 11940 9620 11996
rect 9620 11940 9624 11996
rect 9560 11936 9624 11940
rect 9640 11996 9704 12000
rect 9640 11940 9644 11996
rect 9644 11940 9700 11996
rect 9700 11940 9704 11996
rect 9640 11936 9704 11940
rect 17848 11996 17912 12000
rect 17848 11940 17852 11996
rect 17852 11940 17908 11996
rect 17908 11940 17912 11996
rect 17848 11936 17912 11940
rect 17928 11996 17992 12000
rect 17928 11940 17932 11996
rect 17932 11940 17988 11996
rect 17988 11940 17992 11996
rect 17928 11936 17992 11940
rect 18008 11996 18072 12000
rect 18008 11940 18012 11996
rect 18012 11940 18068 11996
rect 18068 11940 18072 11996
rect 18008 11936 18072 11940
rect 18088 11996 18152 12000
rect 18088 11940 18092 11996
rect 18092 11940 18148 11996
rect 18148 11940 18152 11996
rect 18088 11936 18152 11940
rect 26296 11996 26360 12000
rect 26296 11940 26300 11996
rect 26300 11940 26356 11996
rect 26356 11940 26360 11996
rect 26296 11936 26360 11940
rect 26376 11996 26440 12000
rect 26376 11940 26380 11996
rect 26380 11940 26436 11996
rect 26436 11940 26440 11996
rect 26376 11936 26440 11940
rect 26456 11996 26520 12000
rect 26456 11940 26460 11996
rect 26460 11940 26516 11996
rect 26516 11940 26520 11996
rect 26456 11936 26520 11940
rect 26536 11996 26600 12000
rect 26536 11940 26540 11996
rect 26540 11940 26596 11996
rect 26596 11940 26600 11996
rect 26536 11936 26600 11940
rect 5176 11452 5240 11456
rect 5176 11396 5180 11452
rect 5180 11396 5236 11452
rect 5236 11396 5240 11452
rect 5176 11392 5240 11396
rect 5256 11452 5320 11456
rect 5256 11396 5260 11452
rect 5260 11396 5316 11452
rect 5316 11396 5320 11452
rect 5256 11392 5320 11396
rect 5336 11452 5400 11456
rect 5336 11396 5340 11452
rect 5340 11396 5396 11452
rect 5396 11396 5400 11452
rect 5336 11392 5400 11396
rect 5416 11452 5480 11456
rect 5416 11396 5420 11452
rect 5420 11396 5476 11452
rect 5476 11396 5480 11452
rect 5416 11392 5480 11396
rect 13624 11452 13688 11456
rect 13624 11396 13628 11452
rect 13628 11396 13684 11452
rect 13684 11396 13688 11452
rect 13624 11392 13688 11396
rect 13704 11452 13768 11456
rect 13704 11396 13708 11452
rect 13708 11396 13764 11452
rect 13764 11396 13768 11452
rect 13704 11392 13768 11396
rect 13784 11452 13848 11456
rect 13784 11396 13788 11452
rect 13788 11396 13844 11452
rect 13844 11396 13848 11452
rect 13784 11392 13848 11396
rect 13864 11452 13928 11456
rect 13864 11396 13868 11452
rect 13868 11396 13924 11452
rect 13924 11396 13928 11452
rect 13864 11392 13928 11396
rect 22072 11452 22136 11456
rect 22072 11396 22076 11452
rect 22076 11396 22132 11452
rect 22132 11396 22136 11452
rect 22072 11392 22136 11396
rect 22152 11452 22216 11456
rect 22152 11396 22156 11452
rect 22156 11396 22212 11452
rect 22212 11396 22216 11452
rect 22152 11392 22216 11396
rect 22232 11452 22296 11456
rect 22232 11396 22236 11452
rect 22236 11396 22292 11452
rect 22292 11396 22296 11452
rect 22232 11392 22296 11396
rect 22312 11452 22376 11456
rect 22312 11396 22316 11452
rect 22316 11396 22372 11452
rect 22372 11396 22376 11452
rect 22312 11392 22376 11396
rect 30520 11452 30584 11456
rect 30520 11396 30524 11452
rect 30524 11396 30580 11452
rect 30580 11396 30584 11452
rect 30520 11392 30584 11396
rect 30600 11452 30664 11456
rect 30600 11396 30604 11452
rect 30604 11396 30660 11452
rect 30660 11396 30664 11452
rect 30600 11392 30664 11396
rect 30680 11452 30744 11456
rect 30680 11396 30684 11452
rect 30684 11396 30740 11452
rect 30740 11396 30744 11452
rect 30680 11392 30744 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 9400 10908 9464 10912
rect 9400 10852 9404 10908
rect 9404 10852 9460 10908
rect 9460 10852 9464 10908
rect 9400 10848 9464 10852
rect 9480 10908 9544 10912
rect 9480 10852 9484 10908
rect 9484 10852 9540 10908
rect 9540 10852 9544 10908
rect 9480 10848 9544 10852
rect 9560 10908 9624 10912
rect 9560 10852 9564 10908
rect 9564 10852 9620 10908
rect 9620 10852 9624 10908
rect 9560 10848 9624 10852
rect 9640 10908 9704 10912
rect 9640 10852 9644 10908
rect 9644 10852 9700 10908
rect 9700 10852 9704 10908
rect 9640 10848 9704 10852
rect 17848 10908 17912 10912
rect 17848 10852 17852 10908
rect 17852 10852 17908 10908
rect 17908 10852 17912 10908
rect 17848 10848 17912 10852
rect 17928 10908 17992 10912
rect 17928 10852 17932 10908
rect 17932 10852 17988 10908
rect 17988 10852 17992 10908
rect 17928 10848 17992 10852
rect 18008 10908 18072 10912
rect 18008 10852 18012 10908
rect 18012 10852 18068 10908
rect 18068 10852 18072 10908
rect 18008 10848 18072 10852
rect 18088 10908 18152 10912
rect 18088 10852 18092 10908
rect 18092 10852 18148 10908
rect 18148 10852 18152 10908
rect 18088 10848 18152 10852
rect 26296 10908 26360 10912
rect 26296 10852 26300 10908
rect 26300 10852 26356 10908
rect 26356 10852 26360 10908
rect 26296 10848 26360 10852
rect 26376 10908 26440 10912
rect 26376 10852 26380 10908
rect 26380 10852 26436 10908
rect 26436 10852 26440 10908
rect 26376 10848 26440 10852
rect 26456 10908 26520 10912
rect 26456 10852 26460 10908
rect 26460 10852 26516 10908
rect 26516 10852 26520 10908
rect 26456 10848 26520 10852
rect 26536 10908 26600 10912
rect 26536 10852 26540 10908
rect 26540 10852 26596 10908
rect 26596 10852 26600 10908
rect 26536 10848 26600 10852
rect 5176 10364 5240 10368
rect 5176 10308 5180 10364
rect 5180 10308 5236 10364
rect 5236 10308 5240 10364
rect 5176 10304 5240 10308
rect 5256 10364 5320 10368
rect 5256 10308 5260 10364
rect 5260 10308 5316 10364
rect 5316 10308 5320 10364
rect 5256 10304 5320 10308
rect 5336 10364 5400 10368
rect 5336 10308 5340 10364
rect 5340 10308 5396 10364
rect 5396 10308 5400 10364
rect 5336 10304 5400 10308
rect 5416 10364 5480 10368
rect 5416 10308 5420 10364
rect 5420 10308 5476 10364
rect 5476 10308 5480 10364
rect 5416 10304 5480 10308
rect 13624 10364 13688 10368
rect 13624 10308 13628 10364
rect 13628 10308 13684 10364
rect 13684 10308 13688 10364
rect 13624 10304 13688 10308
rect 13704 10364 13768 10368
rect 13704 10308 13708 10364
rect 13708 10308 13764 10364
rect 13764 10308 13768 10364
rect 13704 10304 13768 10308
rect 13784 10364 13848 10368
rect 13784 10308 13788 10364
rect 13788 10308 13844 10364
rect 13844 10308 13848 10364
rect 13784 10304 13848 10308
rect 13864 10364 13928 10368
rect 13864 10308 13868 10364
rect 13868 10308 13924 10364
rect 13924 10308 13928 10364
rect 13864 10304 13928 10308
rect 22072 10364 22136 10368
rect 22072 10308 22076 10364
rect 22076 10308 22132 10364
rect 22132 10308 22136 10364
rect 22072 10304 22136 10308
rect 22152 10364 22216 10368
rect 22152 10308 22156 10364
rect 22156 10308 22212 10364
rect 22212 10308 22216 10364
rect 22152 10304 22216 10308
rect 22232 10364 22296 10368
rect 22232 10308 22236 10364
rect 22236 10308 22292 10364
rect 22292 10308 22296 10364
rect 22232 10304 22296 10308
rect 22312 10364 22376 10368
rect 22312 10308 22316 10364
rect 22316 10308 22372 10364
rect 22372 10308 22376 10364
rect 22312 10304 22376 10308
rect 30520 10364 30584 10368
rect 30520 10308 30524 10364
rect 30524 10308 30580 10364
rect 30580 10308 30584 10364
rect 30520 10304 30584 10308
rect 30600 10364 30664 10368
rect 30600 10308 30604 10364
rect 30604 10308 30660 10364
rect 30660 10308 30664 10364
rect 30600 10304 30664 10308
rect 30680 10364 30744 10368
rect 30680 10308 30684 10364
rect 30684 10308 30740 10364
rect 30740 10308 30744 10364
rect 30680 10304 30744 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 9400 9820 9464 9824
rect 9400 9764 9404 9820
rect 9404 9764 9460 9820
rect 9460 9764 9464 9820
rect 9400 9760 9464 9764
rect 9480 9820 9544 9824
rect 9480 9764 9484 9820
rect 9484 9764 9540 9820
rect 9540 9764 9544 9820
rect 9480 9760 9544 9764
rect 9560 9820 9624 9824
rect 9560 9764 9564 9820
rect 9564 9764 9620 9820
rect 9620 9764 9624 9820
rect 9560 9760 9624 9764
rect 9640 9820 9704 9824
rect 9640 9764 9644 9820
rect 9644 9764 9700 9820
rect 9700 9764 9704 9820
rect 9640 9760 9704 9764
rect 17848 9820 17912 9824
rect 17848 9764 17852 9820
rect 17852 9764 17908 9820
rect 17908 9764 17912 9820
rect 17848 9760 17912 9764
rect 17928 9820 17992 9824
rect 17928 9764 17932 9820
rect 17932 9764 17988 9820
rect 17988 9764 17992 9820
rect 17928 9760 17992 9764
rect 18008 9820 18072 9824
rect 18008 9764 18012 9820
rect 18012 9764 18068 9820
rect 18068 9764 18072 9820
rect 18008 9760 18072 9764
rect 18088 9820 18152 9824
rect 18088 9764 18092 9820
rect 18092 9764 18148 9820
rect 18148 9764 18152 9820
rect 18088 9760 18152 9764
rect 26296 9820 26360 9824
rect 26296 9764 26300 9820
rect 26300 9764 26356 9820
rect 26356 9764 26360 9820
rect 26296 9760 26360 9764
rect 26376 9820 26440 9824
rect 26376 9764 26380 9820
rect 26380 9764 26436 9820
rect 26436 9764 26440 9820
rect 26376 9760 26440 9764
rect 26456 9820 26520 9824
rect 26456 9764 26460 9820
rect 26460 9764 26516 9820
rect 26516 9764 26520 9820
rect 26456 9760 26520 9764
rect 26536 9820 26600 9824
rect 26536 9764 26540 9820
rect 26540 9764 26596 9820
rect 26596 9764 26600 9820
rect 26536 9760 26600 9764
rect 5176 9276 5240 9280
rect 5176 9220 5180 9276
rect 5180 9220 5236 9276
rect 5236 9220 5240 9276
rect 5176 9216 5240 9220
rect 5256 9276 5320 9280
rect 5256 9220 5260 9276
rect 5260 9220 5316 9276
rect 5316 9220 5320 9276
rect 5256 9216 5320 9220
rect 5336 9276 5400 9280
rect 5336 9220 5340 9276
rect 5340 9220 5396 9276
rect 5396 9220 5400 9276
rect 5336 9216 5400 9220
rect 5416 9276 5480 9280
rect 5416 9220 5420 9276
rect 5420 9220 5476 9276
rect 5476 9220 5480 9276
rect 5416 9216 5480 9220
rect 13624 9276 13688 9280
rect 13624 9220 13628 9276
rect 13628 9220 13684 9276
rect 13684 9220 13688 9276
rect 13624 9216 13688 9220
rect 13704 9276 13768 9280
rect 13704 9220 13708 9276
rect 13708 9220 13764 9276
rect 13764 9220 13768 9276
rect 13704 9216 13768 9220
rect 13784 9276 13848 9280
rect 13784 9220 13788 9276
rect 13788 9220 13844 9276
rect 13844 9220 13848 9276
rect 13784 9216 13848 9220
rect 13864 9276 13928 9280
rect 13864 9220 13868 9276
rect 13868 9220 13924 9276
rect 13924 9220 13928 9276
rect 13864 9216 13928 9220
rect 22072 9276 22136 9280
rect 22072 9220 22076 9276
rect 22076 9220 22132 9276
rect 22132 9220 22136 9276
rect 22072 9216 22136 9220
rect 22152 9276 22216 9280
rect 22152 9220 22156 9276
rect 22156 9220 22212 9276
rect 22212 9220 22216 9276
rect 22152 9216 22216 9220
rect 22232 9276 22296 9280
rect 22232 9220 22236 9276
rect 22236 9220 22292 9276
rect 22292 9220 22296 9276
rect 22232 9216 22296 9220
rect 22312 9276 22376 9280
rect 22312 9220 22316 9276
rect 22316 9220 22372 9276
rect 22372 9220 22376 9276
rect 22312 9216 22376 9220
rect 30520 9276 30584 9280
rect 30520 9220 30524 9276
rect 30524 9220 30580 9276
rect 30580 9220 30584 9276
rect 30520 9216 30584 9220
rect 30600 9276 30664 9280
rect 30600 9220 30604 9276
rect 30604 9220 30660 9276
rect 30660 9220 30664 9276
rect 30600 9216 30664 9220
rect 30680 9276 30744 9280
rect 30680 9220 30684 9276
rect 30684 9220 30740 9276
rect 30740 9220 30744 9276
rect 30680 9216 30744 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 9400 8732 9464 8736
rect 9400 8676 9404 8732
rect 9404 8676 9460 8732
rect 9460 8676 9464 8732
rect 9400 8672 9464 8676
rect 9480 8732 9544 8736
rect 9480 8676 9484 8732
rect 9484 8676 9540 8732
rect 9540 8676 9544 8732
rect 9480 8672 9544 8676
rect 9560 8732 9624 8736
rect 9560 8676 9564 8732
rect 9564 8676 9620 8732
rect 9620 8676 9624 8732
rect 9560 8672 9624 8676
rect 9640 8732 9704 8736
rect 9640 8676 9644 8732
rect 9644 8676 9700 8732
rect 9700 8676 9704 8732
rect 9640 8672 9704 8676
rect 17848 8732 17912 8736
rect 17848 8676 17852 8732
rect 17852 8676 17908 8732
rect 17908 8676 17912 8732
rect 17848 8672 17912 8676
rect 17928 8732 17992 8736
rect 17928 8676 17932 8732
rect 17932 8676 17988 8732
rect 17988 8676 17992 8732
rect 17928 8672 17992 8676
rect 18008 8732 18072 8736
rect 18008 8676 18012 8732
rect 18012 8676 18068 8732
rect 18068 8676 18072 8732
rect 18008 8672 18072 8676
rect 18088 8732 18152 8736
rect 18088 8676 18092 8732
rect 18092 8676 18148 8732
rect 18148 8676 18152 8732
rect 18088 8672 18152 8676
rect 26296 8732 26360 8736
rect 26296 8676 26300 8732
rect 26300 8676 26356 8732
rect 26356 8676 26360 8732
rect 26296 8672 26360 8676
rect 26376 8732 26440 8736
rect 26376 8676 26380 8732
rect 26380 8676 26436 8732
rect 26436 8676 26440 8732
rect 26376 8672 26440 8676
rect 26456 8732 26520 8736
rect 26456 8676 26460 8732
rect 26460 8676 26516 8732
rect 26516 8676 26520 8732
rect 26456 8672 26520 8676
rect 26536 8732 26600 8736
rect 26536 8676 26540 8732
rect 26540 8676 26596 8732
rect 26596 8676 26600 8732
rect 26536 8672 26600 8676
rect 5176 8188 5240 8192
rect 5176 8132 5180 8188
rect 5180 8132 5236 8188
rect 5236 8132 5240 8188
rect 5176 8128 5240 8132
rect 5256 8188 5320 8192
rect 5256 8132 5260 8188
rect 5260 8132 5316 8188
rect 5316 8132 5320 8188
rect 5256 8128 5320 8132
rect 5336 8188 5400 8192
rect 5336 8132 5340 8188
rect 5340 8132 5396 8188
rect 5396 8132 5400 8188
rect 5336 8128 5400 8132
rect 5416 8188 5480 8192
rect 5416 8132 5420 8188
rect 5420 8132 5476 8188
rect 5476 8132 5480 8188
rect 5416 8128 5480 8132
rect 13624 8188 13688 8192
rect 13624 8132 13628 8188
rect 13628 8132 13684 8188
rect 13684 8132 13688 8188
rect 13624 8128 13688 8132
rect 13704 8188 13768 8192
rect 13704 8132 13708 8188
rect 13708 8132 13764 8188
rect 13764 8132 13768 8188
rect 13704 8128 13768 8132
rect 13784 8188 13848 8192
rect 13784 8132 13788 8188
rect 13788 8132 13844 8188
rect 13844 8132 13848 8188
rect 13784 8128 13848 8132
rect 13864 8188 13928 8192
rect 13864 8132 13868 8188
rect 13868 8132 13924 8188
rect 13924 8132 13928 8188
rect 13864 8128 13928 8132
rect 22072 8188 22136 8192
rect 22072 8132 22076 8188
rect 22076 8132 22132 8188
rect 22132 8132 22136 8188
rect 22072 8128 22136 8132
rect 22152 8188 22216 8192
rect 22152 8132 22156 8188
rect 22156 8132 22212 8188
rect 22212 8132 22216 8188
rect 22152 8128 22216 8132
rect 22232 8188 22296 8192
rect 22232 8132 22236 8188
rect 22236 8132 22292 8188
rect 22292 8132 22296 8188
rect 22232 8128 22296 8132
rect 22312 8188 22376 8192
rect 22312 8132 22316 8188
rect 22316 8132 22372 8188
rect 22372 8132 22376 8188
rect 22312 8128 22376 8132
rect 30520 8188 30584 8192
rect 30520 8132 30524 8188
rect 30524 8132 30580 8188
rect 30580 8132 30584 8188
rect 30520 8128 30584 8132
rect 30600 8188 30664 8192
rect 30600 8132 30604 8188
rect 30604 8132 30660 8188
rect 30660 8132 30664 8188
rect 30600 8128 30664 8132
rect 30680 8188 30744 8192
rect 30680 8132 30684 8188
rect 30684 8132 30740 8188
rect 30740 8132 30744 8188
rect 30680 8128 30744 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 9400 7644 9464 7648
rect 9400 7588 9404 7644
rect 9404 7588 9460 7644
rect 9460 7588 9464 7644
rect 9400 7584 9464 7588
rect 9480 7644 9544 7648
rect 9480 7588 9484 7644
rect 9484 7588 9540 7644
rect 9540 7588 9544 7644
rect 9480 7584 9544 7588
rect 9560 7644 9624 7648
rect 9560 7588 9564 7644
rect 9564 7588 9620 7644
rect 9620 7588 9624 7644
rect 9560 7584 9624 7588
rect 9640 7644 9704 7648
rect 9640 7588 9644 7644
rect 9644 7588 9700 7644
rect 9700 7588 9704 7644
rect 9640 7584 9704 7588
rect 17848 7644 17912 7648
rect 17848 7588 17852 7644
rect 17852 7588 17908 7644
rect 17908 7588 17912 7644
rect 17848 7584 17912 7588
rect 17928 7644 17992 7648
rect 17928 7588 17932 7644
rect 17932 7588 17988 7644
rect 17988 7588 17992 7644
rect 17928 7584 17992 7588
rect 18008 7644 18072 7648
rect 18008 7588 18012 7644
rect 18012 7588 18068 7644
rect 18068 7588 18072 7644
rect 18008 7584 18072 7588
rect 18088 7644 18152 7648
rect 18088 7588 18092 7644
rect 18092 7588 18148 7644
rect 18148 7588 18152 7644
rect 18088 7584 18152 7588
rect 26296 7644 26360 7648
rect 26296 7588 26300 7644
rect 26300 7588 26356 7644
rect 26356 7588 26360 7644
rect 26296 7584 26360 7588
rect 26376 7644 26440 7648
rect 26376 7588 26380 7644
rect 26380 7588 26436 7644
rect 26436 7588 26440 7644
rect 26376 7584 26440 7588
rect 26456 7644 26520 7648
rect 26456 7588 26460 7644
rect 26460 7588 26516 7644
rect 26516 7588 26520 7644
rect 26456 7584 26520 7588
rect 26536 7644 26600 7648
rect 26536 7588 26540 7644
rect 26540 7588 26596 7644
rect 26596 7588 26600 7644
rect 26536 7584 26600 7588
rect 5176 7100 5240 7104
rect 5176 7044 5180 7100
rect 5180 7044 5236 7100
rect 5236 7044 5240 7100
rect 5176 7040 5240 7044
rect 5256 7100 5320 7104
rect 5256 7044 5260 7100
rect 5260 7044 5316 7100
rect 5316 7044 5320 7100
rect 5256 7040 5320 7044
rect 5336 7100 5400 7104
rect 5336 7044 5340 7100
rect 5340 7044 5396 7100
rect 5396 7044 5400 7100
rect 5336 7040 5400 7044
rect 5416 7100 5480 7104
rect 5416 7044 5420 7100
rect 5420 7044 5476 7100
rect 5476 7044 5480 7100
rect 5416 7040 5480 7044
rect 13624 7100 13688 7104
rect 13624 7044 13628 7100
rect 13628 7044 13684 7100
rect 13684 7044 13688 7100
rect 13624 7040 13688 7044
rect 13704 7100 13768 7104
rect 13704 7044 13708 7100
rect 13708 7044 13764 7100
rect 13764 7044 13768 7100
rect 13704 7040 13768 7044
rect 13784 7100 13848 7104
rect 13784 7044 13788 7100
rect 13788 7044 13844 7100
rect 13844 7044 13848 7100
rect 13784 7040 13848 7044
rect 13864 7100 13928 7104
rect 13864 7044 13868 7100
rect 13868 7044 13924 7100
rect 13924 7044 13928 7100
rect 13864 7040 13928 7044
rect 22072 7100 22136 7104
rect 22072 7044 22076 7100
rect 22076 7044 22132 7100
rect 22132 7044 22136 7100
rect 22072 7040 22136 7044
rect 22152 7100 22216 7104
rect 22152 7044 22156 7100
rect 22156 7044 22212 7100
rect 22212 7044 22216 7100
rect 22152 7040 22216 7044
rect 22232 7100 22296 7104
rect 22232 7044 22236 7100
rect 22236 7044 22292 7100
rect 22292 7044 22296 7100
rect 22232 7040 22296 7044
rect 22312 7100 22376 7104
rect 22312 7044 22316 7100
rect 22316 7044 22372 7100
rect 22372 7044 22376 7100
rect 22312 7040 22376 7044
rect 30520 7100 30584 7104
rect 30520 7044 30524 7100
rect 30524 7044 30580 7100
rect 30580 7044 30584 7100
rect 30520 7040 30584 7044
rect 30600 7100 30664 7104
rect 30600 7044 30604 7100
rect 30604 7044 30660 7100
rect 30660 7044 30664 7100
rect 30600 7040 30664 7044
rect 30680 7100 30744 7104
rect 30680 7044 30684 7100
rect 30684 7044 30740 7100
rect 30740 7044 30744 7100
rect 30680 7040 30744 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 9400 6556 9464 6560
rect 9400 6500 9404 6556
rect 9404 6500 9460 6556
rect 9460 6500 9464 6556
rect 9400 6496 9464 6500
rect 9480 6556 9544 6560
rect 9480 6500 9484 6556
rect 9484 6500 9540 6556
rect 9540 6500 9544 6556
rect 9480 6496 9544 6500
rect 9560 6556 9624 6560
rect 9560 6500 9564 6556
rect 9564 6500 9620 6556
rect 9620 6500 9624 6556
rect 9560 6496 9624 6500
rect 9640 6556 9704 6560
rect 9640 6500 9644 6556
rect 9644 6500 9700 6556
rect 9700 6500 9704 6556
rect 9640 6496 9704 6500
rect 17848 6556 17912 6560
rect 17848 6500 17852 6556
rect 17852 6500 17908 6556
rect 17908 6500 17912 6556
rect 17848 6496 17912 6500
rect 17928 6556 17992 6560
rect 17928 6500 17932 6556
rect 17932 6500 17988 6556
rect 17988 6500 17992 6556
rect 17928 6496 17992 6500
rect 18008 6556 18072 6560
rect 18008 6500 18012 6556
rect 18012 6500 18068 6556
rect 18068 6500 18072 6556
rect 18008 6496 18072 6500
rect 18088 6556 18152 6560
rect 18088 6500 18092 6556
rect 18092 6500 18148 6556
rect 18148 6500 18152 6556
rect 18088 6496 18152 6500
rect 26296 6556 26360 6560
rect 26296 6500 26300 6556
rect 26300 6500 26356 6556
rect 26356 6500 26360 6556
rect 26296 6496 26360 6500
rect 26376 6556 26440 6560
rect 26376 6500 26380 6556
rect 26380 6500 26436 6556
rect 26436 6500 26440 6556
rect 26376 6496 26440 6500
rect 26456 6556 26520 6560
rect 26456 6500 26460 6556
rect 26460 6500 26516 6556
rect 26516 6500 26520 6556
rect 26456 6496 26520 6500
rect 26536 6556 26600 6560
rect 26536 6500 26540 6556
rect 26540 6500 26596 6556
rect 26596 6500 26600 6556
rect 26536 6496 26600 6500
rect 5176 6012 5240 6016
rect 5176 5956 5180 6012
rect 5180 5956 5236 6012
rect 5236 5956 5240 6012
rect 5176 5952 5240 5956
rect 5256 6012 5320 6016
rect 5256 5956 5260 6012
rect 5260 5956 5316 6012
rect 5316 5956 5320 6012
rect 5256 5952 5320 5956
rect 5336 6012 5400 6016
rect 5336 5956 5340 6012
rect 5340 5956 5396 6012
rect 5396 5956 5400 6012
rect 5336 5952 5400 5956
rect 5416 6012 5480 6016
rect 5416 5956 5420 6012
rect 5420 5956 5476 6012
rect 5476 5956 5480 6012
rect 5416 5952 5480 5956
rect 13624 6012 13688 6016
rect 13624 5956 13628 6012
rect 13628 5956 13684 6012
rect 13684 5956 13688 6012
rect 13624 5952 13688 5956
rect 13704 6012 13768 6016
rect 13704 5956 13708 6012
rect 13708 5956 13764 6012
rect 13764 5956 13768 6012
rect 13704 5952 13768 5956
rect 13784 6012 13848 6016
rect 13784 5956 13788 6012
rect 13788 5956 13844 6012
rect 13844 5956 13848 6012
rect 13784 5952 13848 5956
rect 13864 6012 13928 6016
rect 13864 5956 13868 6012
rect 13868 5956 13924 6012
rect 13924 5956 13928 6012
rect 13864 5952 13928 5956
rect 22072 6012 22136 6016
rect 22072 5956 22076 6012
rect 22076 5956 22132 6012
rect 22132 5956 22136 6012
rect 22072 5952 22136 5956
rect 22152 6012 22216 6016
rect 22152 5956 22156 6012
rect 22156 5956 22212 6012
rect 22212 5956 22216 6012
rect 22152 5952 22216 5956
rect 22232 6012 22296 6016
rect 22232 5956 22236 6012
rect 22236 5956 22292 6012
rect 22292 5956 22296 6012
rect 22232 5952 22296 5956
rect 22312 6012 22376 6016
rect 22312 5956 22316 6012
rect 22316 5956 22372 6012
rect 22372 5956 22376 6012
rect 22312 5952 22376 5956
rect 30520 6012 30584 6016
rect 30520 5956 30524 6012
rect 30524 5956 30580 6012
rect 30580 5956 30584 6012
rect 30520 5952 30584 5956
rect 30600 6012 30664 6016
rect 30600 5956 30604 6012
rect 30604 5956 30660 6012
rect 30660 5956 30664 6012
rect 30600 5952 30664 5956
rect 30680 6012 30744 6016
rect 30680 5956 30684 6012
rect 30684 5956 30740 6012
rect 30740 5956 30744 6012
rect 30680 5952 30744 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 9400 5468 9464 5472
rect 9400 5412 9404 5468
rect 9404 5412 9460 5468
rect 9460 5412 9464 5468
rect 9400 5408 9464 5412
rect 9480 5468 9544 5472
rect 9480 5412 9484 5468
rect 9484 5412 9540 5468
rect 9540 5412 9544 5468
rect 9480 5408 9544 5412
rect 9560 5468 9624 5472
rect 9560 5412 9564 5468
rect 9564 5412 9620 5468
rect 9620 5412 9624 5468
rect 9560 5408 9624 5412
rect 9640 5468 9704 5472
rect 9640 5412 9644 5468
rect 9644 5412 9700 5468
rect 9700 5412 9704 5468
rect 9640 5408 9704 5412
rect 17848 5468 17912 5472
rect 17848 5412 17852 5468
rect 17852 5412 17908 5468
rect 17908 5412 17912 5468
rect 17848 5408 17912 5412
rect 17928 5468 17992 5472
rect 17928 5412 17932 5468
rect 17932 5412 17988 5468
rect 17988 5412 17992 5468
rect 17928 5408 17992 5412
rect 18008 5468 18072 5472
rect 18008 5412 18012 5468
rect 18012 5412 18068 5468
rect 18068 5412 18072 5468
rect 18008 5408 18072 5412
rect 18088 5468 18152 5472
rect 18088 5412 18092 5468
rect 18092 5412 18148 5468
rect 18148 5412 18152 5468
rect 18088 5408 18152 5412
rect 26296 5468 26360 5472
rect 26296 5412 26300 5468
rect 26300 5412 26356 5468
rect 26356 5412 26360 5468
rect 26296 5408 26360 5412
rect 26376 5468 26440 5472
rect 26376 5412 26380 5468
rect 26380 5412 26436 5468
rect 26436 5412 26440 5468
rect 26376 5408 26440 5412
rect 26456 5468 26520 5472
rect 26456 5412 26460 5468
rect 26460 5412 26516 5468
rect 26516 5412 26520 5468
rect 26456 5408 26520 5412
rect 26536 5468 26600 5472
rect 26536 5412 26540 5468
rect 26540 5412 26596 5468
rect 26596 5412 26600 5468
rect 26536 5408 26600 5412
rect 5176 4924 5240 4928
rect 5176 4868 5180 4924
rect 5180 4868 5236 4924
rect 5236 4868 5240 4924
rect 5176 4864 5240 4868
rect 5256 4924 5320 4928
rect 5256 4868 5260 4924
rect 5260 4868 5316 4924
rect 5316 4868 5320 4924
rect 5256 4864 5320 4868
rect 5336 4924 5400 4928
rect 5336 4868 5340 4924
rect 5340 4868 5396 4924
rect 5396 4868 5400 4924
rect 5336 4864 5400 4868
rect 5416 4924 5480 4928
rect 5416 4868 5420 4924
rect 5420 4868 5476 4924
rect 5476 4868 5480 4924
rect 5416 4864 5480 4868
rect 13624 4924 13688 4928
rect 13624 4868 13628 4924
rect 13628 4868 13684 4924
rect 13684 4868 13688 4924
rect 13624 4864 13688 4868
rect 13704 4924 13768 4928
rect 13704 4868 13708 4924
rect 13708 4868 13764 4924
rect 13764 4868 13768 4924
rect 13704 4864 13768 4868
rect 13784 4924 13848 4928
rect 13784 4868 13788 4924
rect 13788 4868 13844 4924
rect 13844 4868 13848 4924
rect 13784 4864 13848 4868
rect 13864 4924 13928 4928
rect 13864 4868 13868 4924
rect 13868 4868 13924 4924
rect 13924 4868 13928 4924
rect 13864 4864 13928 4868
rect 22072 4924 22136 4928
rect 22072 4868 22076 4924
rect 22076 4868 22132 4924
rect 22132 4868 22136 4924
rect 22072 4864 22136 4868
rect 22152 4924 22216 4928
rect 22152 4868 22156 4924
rect 22156 4868 22212 4924
rect 22212 4868 22216 4924
rect 22152 4864 22216 4868
rect 22232 4924 22296 4928
rect 22232 4868 22236 4924
rect 22236 4868 22292 4924
rect 22292 4868 22296 4924
rect 22232 4864 22296 4868
rect 22312 4924 22376 4928
rect 22312 4868 22316 4924
rect 22316 4868 22372 4924
rect 22372 4868 22376 4924
rect 22312 4864 22376 4868
rect 30520 4924 30584 4928
rect 30520 4868 30524 4924
rect 30524 4868 30580 4924
rect 30580 4868 30584 4924
rect 30520 4864 30584 4868
rect 30600 4924 30664 4928
rect 30600 4868 30604 4924
rect 30604 4868 30660 4924
rect 30660 4868 30664 4924
rect 30600 4864 30664 4868
rect 30680 4924 30744 4928
rect 30680 4868 30684 4924
rect 30684 4868 30740 4924
rect 30740 4868 30744 4924
rect 30680 4864 30744 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 9400 4380 9464 4384
rect 9400 4324 9404 4380
rect 9404 4324 9460 4380
rect 9460 4324 9464 4380
rect 9400 4320 9464 4324
rect 9480 4380 9544 4384
rect 9480 4324 9484 4380
rect 9484 4324 9540 4380
rect 9540 4324 9544 4380
rect 9480 4320 9544 4324
rect 9560 4380 9624 4384
rect 9560 4324 9564 4380
rect 9564 4324 9620 4380
rect 9620 4324 9624 4380
rect 9560 4320 9624 4324
rect 9640 4380 9704 4384
rect 9640 4324 9644 4380
rect 9644 4324 9700 4380
rect 9700 4324 9704 4380
rect 9640 4320 9704 4324
rect 17848 4380 17912 4384
rect 17848 4324 17852 4380
rect 17852 4324 17908 4380
rect 17908 4324 17912 4380
rect 17848 4320 17912 4324
rect 17928 4380 17992 4384
rect 17928 4324 17932 4380
rect 17932 4324 17988 4380
rect 17988 4324 17992 4380
rect 17928 4320 17992 4324
rect 18008 4380 18072 4384
rect 18008 4324 18012 4380
rect 18012 4324 18068 4380
rect 18068 4324 18072 4380
rect 18008 4320 18072 4324
rect 18088 4380 18152 4384
rect 18088 4324 18092 4380
rect 18092 4324 18148 4380
rect 18148 4324 18152 4380
rect 18088 4320 18152 4324
rect 26296 4380 26360 4384
rect 26296 4324 26300 4380
rect 26300 4324 26356 4380
rect 26356 4324 26360 4380
rect 26296 4320 26360 4324
rect 26376 4380 26440 4384
rect 26376 4324 26380 4380
rect 26380 4324 26436 4380
rect 26436 4324 26440 4380
rect 26376 4320 26440 4324
rect 26456 4380 26520 4384
rect 26456 4324 26460 4380
rect 26460 4324 26516 4380
rect 26516 4324 26520 4380
rect 26456 4320 26520 4324
rect 26536 4380 26600 4384
rect 26536 4324 26540 4380
rect 26540 4324 26596 4380
rect 26596 4324 26600 4380
rect 26536 4320 26600 4324
rect 5176 3836 5240 3840
rect 5176 3780 5180 3836
rect 5180 3780 5236 3836
rect 5236 3780 5240 3836
rect 5176 3776 5240 3780
rect 5256 3836 5320 3840
rect 5256 3780 5260 3836
rect 5260 3780 5316 3836
rect 5316 3780 5320 3836
rect 5256 3776 5320 3780
rect 5336 3836 5400 3840
rect 5336 3780 5340 3836
rect 5340 3780 5396 3836
rect 5396 3780 5400 3836
rect 5336 3776 5400 3780
rect 5416 3836 5480 3840
rect 5416 3780 5420 3836
rect 5420 3780 5476 3836
rect 5476 3780 5480 3836
rect 5416 3776 5480 3780
rect 13624 3836 13688 3840
rect 13624 3780 13628 3836
rect 13628 3780 13684 3836
rect 13684 3780 13688 3836
rect 13624 3776 13688 3780
rect 13704 3836 13768 3840
rect 13704 3780 13708 3836
rect 13708 3780 13764 3836
rect 13764 3780 13768 3836
rect 13704 3776 13768 3780
rect 13784 3836 13848 3840
rect 13784 3780 13788 3836
rect 13788 3780 13844 3836
rect 13844 3780 13848 3836
rect 13784 3776 13848 3780
rect 13864 3836 13928 3840
rect 13864 3780 13868 3836
rect 13868 3780 13924 3836
rect 13924 3780 13928 3836
rect 13864 3776 13928 3780
rect 22072 3836 22136 3840
rect 22072 3780 22076 3836
rect 22076 3780 22132 3836
rect 22132 3780 22136 3836
rect 22072 3776 22136 3780
rect 22152 3836 22216 3840
rect 22152 3780 22156 3836
rect 22156 3780 22212 3836
rect 22212 3780 22216 3836
rect 22152 3776 22216 3780
rect 22232 3836 22296 3840
rect 22232 3780 22236 3836
rect 22236 3780 22292 3836
rect 22292 3780 22296 3836
rect 22232 3776 22296 3780
rect 22312 3836 22376 3840
rect 22312 3780 22316 3836
rect 22316 3780 22372 3836
rect 22372 3780 22376 3836
rect 22312 3776 22376 3780
rect 30520 3836 30584 3840
rect 30520 3780 30524 3836
rect 30524 3780 30580 3836
rect 30580 3780 30584 3836
rect 30520 3776 30584 3780
rect 30600 3836 30664 3840
rect 30600 3780 30604 3836
rect 30604 3780 30660 3836
rect 30660 3780 30664 3836
rect 30600 3776 30664 3780
rect 30680 3836 30744 3840
rect 30680 3780 30684 3836
rect 30684 3780 30740 3836
rect 30740 3780 30744 3836
rect 30680 3776 30744 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 9400 3292 9464 3296
rect 9400 3236 9404 3292
rect 9404 3236 9460 3292
rect 9460 3236 9464 3292
rect 9400 3232 9464 3236
rect 9480 3292 9544 3296
rect 9480 3236 9484 3292
rect 9484 3236 9540 3292
rect 9540 3236 9544 3292
rect 9480 3232 9544 3236
rect 9560 3292 9624 3296
rect 9560 3236 9564 3292
rect 9564 3236 9620 3292
rect 9620 3236 9624 3292
rect 9560 3232 9624 3236
rect 9640 3292 9704 3296
rect 9640 3236 9644 3292
rect 9644 3236 9700 3292
rect 9700 3236 9704 3292
rect 9640 3232 9704 3236
rect 17848 3292 17912 3296
rect 17848 3236 17852 3292
rect 17852 3236 17908 3292
rect 17908 3236 17912 3292
rect 17848 3232 17912 3236
rect 17928 3292 17992 3296
rect 17928 3236 17932 3292
rect 17932 3236 17988 3292
rect 17988 3236 17992 3292
rect 17928 3232 17992 3236
rect 18008 3292 18072 3296
rect 18008 3236 18012 3292
rect 18012 3236 18068 3292
rect 18068 3236 18072 3292
rect 18008 3232 18072 3236
rect 18088 3292 18152 3296
rect 18088 3236 18092 3292
rect 18092 3236 18148 3292
rect 18148 3236 18152 3292
rect 18088 3232 18152 3236
rect 26296 3292 26360 3296
rect 26296 3236 26300 3292
rect 26300 3236 26356 3292
rect 26356 3236 26360 3292
rect 26296 3232 26360 3236
rect 26376 3292 26440 3296
rect 26376 3236 26380 3292
rect 26380 3236 26436 3292
rect 26436 3236 26440 3292
rect 26376 3232 26440 3236
rect 26456 3292 26520 3296
rect 26456 3236 26460 3292
rect 26460 3236 26516 3292
rect 26516 3236 26520 3292
rect 26456 3232 26520 3236
rect 26536 3292 26600 3296
rect 26536 3236 26540 3292
rect 26540 3236 26596 3292
rect 26596 3236 26600 3292
rect 26536 3232 26600 3236
rect 5176 2748 5240 2752
rect 5176 2692 5180 2748
rect 5180 2692 5236 2748
rect 5236 2692 5240 2748
rect 5176 2688 5240 2692
rect 5256 2748 5320 2752
rect 5256 2692 5260 2748
rect 5260 2692 5316 2748
rect 5316 2692 5320 2748
rect 5256 2688 5320 2692
rect 5336 2748 5400 2752
rect 5336 2692 5340 2748
rect 5340 2692 5396 2748
rect 5396 2692 5400 2748
rect 5336 2688 5400 2692
rect 5416 2748 5480 2752
rect 5416 2692 5420 2748
rect 5420 2692 5476 2748
rect 5476 2692 5480 2748
rect 5416 2688 5480 2692
rect 13624 2748 13688 2752
rect 13624 2692 13628 2748
rect 13628 2692 13684 2748
rect 13684 2692 13688 2748
rect 13624 2688 13688 2692
rect 13704 2748 13768 2752
rect 13704 2692 13708 2748
rect 13708 2692 13764 2748
rect 13764 2692 13768 2748
rect 13704 2688 13768 2692
rect 13784 2748 13848 2752
rect 13784 2692 13788 2748
rect 13788 2692 13844 2748
rect 13844 2692 13848 2748
rect 13784 2688 13848 2692
rect 13864 2748 13928 2752
rect 13864 2692 13868 2748
rect 13868 2692 13924 2748
rect 13924 2692 13928 2748
rect 13864 2688 13928 2692
rect 22072 2748 22136 2752
rect 22072 2692 22076 2748
rect 22076 2692 22132 2748
rect 22132 2692 22136 2748
rect 22072 2688 22136 2692
rect 22152 2748 22216 2752
rect 22152 2692 22156 2748
rect 22156 2692 22212 2748
rect 22212 2692 22216 2748
rect 22152 2688 22216 2692
rect 22232 2748 22296 2752
rect 22232 2692 22236 2748
rect 22236 2692 22292 2748
rect 22292 2692 22296 2748
rect 22232 2688 22296 2692
rect 22312 2748 22376 2752
rect 22312 2692 22316 2748
rect 22316 2692 22372 2748
rect 22372 2692 22376 2748
rect 22312 2688 22376 2692
rect 30520 2748 30584 2752
rect 30520 2692 30524 2748
rect 30524 2692 30580 2748
rect 30580 2692 30584 2748
rect 30520 2688 30584 2692
rect 30600 2748 30664 2752
rect 30600 2692 30604 2748
rect 30604 2692 30660 2748
rect 30660 2692 30664 2748
rect 30600 2688 30664 2692
rect 30680 2748 30744 2752
rect 30680 2692 30684 2748
rect 30684 2692 30740 2748
rect 30740 2692 30744 2748
rect 30680 2688 30744 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 9400 2204 9464 2208
rect 9400 2148 9404 2204
rect 9404 2148 9460 2204
rect 9460 2148 9464 2204
rect 9400 2144 9464 2148
rect 9480 2204 9544 2208
rect 9480 2148 9484 2204
rect 9484 2148 9540 2204
rect 9540 2148 9544 2204
rect 9480 2144 9544 2148
rect 9560 2204 9624 2208
rect 9560 2148 9564 2204
rect 9564 2148 9620 2204
rect 9620 2148 9624 2204
rect 9560 2144 9624 2148
rect 9640 2204 9704 2208
rect 9640 2148 9644 2204
rect 9644 2148 9700 2204
rect 9700 2148 9704 2204
rect 9640 2144 9704 2148
rect 17848 2204 17912 2208
rect 17848 2148 17852 2204
rect 17852 2148 17908 2204
rect 17908 2148 17912 2204
rect 17848 2144 17912 2148
rect 17928 2204 17992 2208
rect 17928 2148 17932 2204
rect 17932 2148 17988 2204
rect 17988 2148 17992 2204
rect 17928 2144 17992 2148
rect 18008 2204 18072 2208
rect 18008 2148 18012 2204
rect 18012 2148 18068 2204
rect 18068 2148 18072 2204
rect 18008 2144 18072 2148
rect 18088 2204 18152 2208
rect 18088 2148 18092 2204
rect 18092 2148 18148 2204
rect 18148 2148 18152 2204
rect 18088 2144 18152 2148
rect 26296 2204 26360 2208
rect 26296 2148 26300 2204
rect 26300 2148 26356 2204
rect 26356 2148 26360 2204
rect 26296 2144 26360 2148
rect 26376 2204 26440 2208
rect 26376 2148 26380 2204
rect 26380 2148 26436 2204
rect 26436 2148 26440 2204
rect 26376 2144 26440 2148
rect 26456 2204 26520 2208
rect 26456 2148 26460 2204
rect 26460 2148 26516 2204
rect 26516 2148 26520 2204
rect 26456 2144 26520 2148
rect 26536 2204 26600 2208
rect 26536 2148 26540 2204
rect 26540 2148 26596 2204
rect 26596 2148 26600 2204
rect 26536 2144 26600 2148
<< metal4 >>
rect 5168 39744 5488 39760
rect 5168 39680 5176 39744
rect 5240 39680 5256 39744
rect 5320 39680 5336 39744
rect 5400 39680 5416 39744
rect 5480 39680 5488 39744
rect 5168 38656 5488 39680
rect 5168 38592 5176 38656
rect 5240 38592 5256 38656
rect 5320 38592 5336 38656
rect 5400 38592 5416 38656
rect 5480 38592 5488 38656
rect 5168 37568 5488 38592
rect 5168 37504 5176 37568
rect 5240 37504 5256 37568
rect 5320 37504 5336 37568
rect 5400 37504 5416 37568
rect 5480 37504 5488 37568
rect 5168 36480 5488 37504
rect 5168 36416 5176 36480
rect 5240 36416 5256 36480
rect 5320 36416 5336 36480
rect 5400 36416 5416 36480
rect 5480 36416 5488 36480
rect 5168 35392 5488 36416
rect 5168 35328 5176 35392
rect 5240 35328 5256 35392
rect 5320 35328 5336 35392
rect 5400 35328 5416 35392
rect 5480 35328 5488 35392
rect 5168 34304 5488 35328
rect 5168 34240 5176 34304
rect 5240 34240 5256 34304
rect 5320 34240 5336 34304
rect 5400 34240 5416 34304
rect 5480 34240 5488 34304
rect 5168 33216 5488 34240
rect 5168 33152 5176 33216
rect 5240 33152 5256 33216
rect 5320 33152 5336 33216
rect 5400 33152 5416 33216
rect 5480 33152 5488 33216
rect 5168 32128 5488 33152
rect 5168 32064 5176 32128
rect 5240 32064 5256 32128
rect 5320 32064 5336 32128
rect 5400 32064 5416 32128
rect 5480 32064 5488 32128
rect 5168 31040 5488 32064
rect 5168 30976 5176 31040
rect 5240 30976 5256 31040
rect 5320 30976 5336 31040
rect 5400 30976 5416 31040
rect 5480 30976 5488 31040
rect 5168 29952 5488 30976
rect 5168 29888 5176 29952
rect 5240 29888 5256 29952
rect 5320 29888 5336 29952
rect 5400 29888 5416 29952
rect 5480 29888 5488 29952
rect 5168 28864 5488 29888
rect 5168 28800 5176 28864
rect 5240 28800 5256 28864
rect 5320 28800 5336 28864
rect 5400 28800 5416 28864
rect 5480 28800 5488 28864
rect 5168 27776 5488 28800
rect 5168 27712 5176 27776
rect 5240 27712 5256 27776
rect 5320 27712 5336 27776
rect 5400 27712 5416 27776
rect 5480 27712 5488 27776
rect 5168 26688 5488 27712
rect 5168 26624 5176 26688
rect 5240 26624 5256 26688
rect 5320 26624 5336 26688
rect 5400 26624 5416 26688
rect 5480 26624 5488 26688
rect 5168 25600 5488 26624
rect 5168 25536 5176 25600
rect 5240 25536 5256 25600
rect 5320 25536 5336 25600
rect 5400 25536 5416 25600
rect 5480 25536 5488 25600
rect 5168 24512 5488 25536
rect 5168 24448 5176 24512
rect 5240 24448 5256 24512
rect 5320 24448 5336 24512
rect 5400 24448 5416 24512
rect 5480 24448 5488 24512
rect 5168 23424 5488 24448
rect 5168 23360 5176 23424
rect 5240 23360 5256 23424
rect 5320 23360 5336 23424
rect 5400 23360 5416 23424
rect 5480 23360 5488 23424
rect 5168 22336 5488 23360
rect 5168 22272 5176 22336
rect 5240 22272 5256 22336
rect 5320 22272 5336 22336
rect 5400 22272 5416 22336
rect 5480 22272 5488 22336
rect 5168 21248 5488 22272
rect 5168 21184 5176 21248
rect 5240 21184 5256 21248
rect 5320 21184 5336 21248
rect 5400 21184 5416 21248
rect 5480 21184 5488 21248
rect 5168 20160 5488 21184
rect 5168 20096 5176 20160
rect 5240 20096 5256 20160
rect 5320 20096 5336 20160
rect 5400 20096 5416 20160
rect 5480 20096 5488 20160
rect 5168 19072 5488 20096
rect 5168 19008 5176 19072
rect 5240 19008 5256 19072
rect 5320 19008 5336 19072
rect 5400 19008 5416 19072
rect 5480 19008 5488 19072
rect 5168 17984 5488 19008
rect 5168 17920 5176 17984
rect 5240 17920 5256 17984
rect 5320 17920 5336 17984
rect 5400 17920 5416 17984
rect 5480 17920 5488 17984
rect 5168 16896 5488 17920
rect 5168 16832 5176 16896
rect 5240 16832 5256 16896
rect 5320 16832 5336 16896
rect 5400 16832 5416 16896
rect 5480 16832 5488 16896
rect 5168 15808 5488 16832
rect 5168 15744 5176 15808
rect 5240 15744 5256 15808
rect 5320 15744 5336 15808
rect 5400 15744 5416 15808
rect 5480 15744 5488 15808
rect 5168 14720 5488 15744
rect 5168 14656 5176 14720
rect 5240 14656 5256 14720
rect 5320 14656 5336 14720
rect 5400 14656 5416 14720
rect 5480 14656 5488 14720
rect 5168 13632 5488 14656
rect 5168 13568 5176 13632
rect 5240 13568 5256 13632
rect 5320 13568 5336 13632
rect 5400 13568 5416 13632
rect 5480 13568 5488 13632
rect 5168 12544 5488 13568
rect 5168 12480 5176 12544
rect 5240 12480 5256 12544
rect 5320 12480 5336 12544
rect 5400 12480 5416 12544
rect 5480 12480 5488 12544
rect 5168 11456 5488 12480
rect 5168 11392 5176 11456
rect 5240 11392 5256 11456
rect 5320 11392 5336 11456
rect 5400 11392 5416 11456
rect 5480 11392 5488 11456
rect 5168 10368 5488 11392
rect 5168 10304 5176 10368
rect 5240 10304 5256 10368
rect 5320 10304 5336 10368
rect 5400 10304 5416 10368
rect 5480 10304 5488 10368
rect 5168 9280 5488 10304
rect 5168 9216 5176 9280
rect 5240 9216 5256 9280
rect 5320 9216 5336 9280
rect 5400 9216 5416 9280
rect 5480 9216 5488 9280
rect 5168 8192 5488 9216
rect 5168 8128 5176 8192
rect 5240 8128 5256 8192
rect 5320 8128 5336 8192
rect 5400 8128 5416 8192
rect 5480 8128 5488 8192
rect 5168 7104 5488 8128
rect 5168 7040 5176 7104
rect 5240 7040 5256 7104
rect 5320 7040 5336 7104
rect 5400 7040 5416 7104
rect 5480 7040 5488 7104
rect 5168 6016 5488 7040
rect 5168 5952 5176 6016
rect 5240 5952 5256 6016
rect 5320 5952 5336 6016
rect 5400 5952 5416 6016
rect 5480 5952 5488 6016
rect 5168 4928 5488 5952
rect 5168 4864 5176 4928
rect 5240 4864 5256 4928
rect 5320 4864 5336 4928
rect 5400 4864 5416 4928
rect 5480 4864 5488 4928
rect 5168 3840 5488 4864
rect 5168 3776 5176 3840
rect 5240 3776 5256 3840
rect 5320 3776 5336 3840
rect 5400 3776 5416 3840
rect 5480 3776 5488 3840
rect 5168 2752 5488 3776
rect 5168 2688 5176 2752
rect 5240 2688 5256 2752
rect 5320 2688 5336 2752
rect 5400 2688 5416 2752
rect 5480 2688 5488 2752
rect 5168 2128 5488 2688
rect 9392 39200 9712 39760
rect 9392 39136 9400 39200
rect 9464 39136 9480 39200
rect 9544 39136 9560 39200
rect 9624 39136 9640 39200
rect 9704 39136 9712 39200
rect 9392 38112 9712 39136
rect 9392 38048 9400 38112
rect 9464 38048 9480 38112
rect 9544 38048 9560 38112
rect 9624 38048 9640 38112
rect 9704 38048 9712 38112
rect 9392 37024 9712 38048
rect 9392 36960 9400 37024
rect 9464 36960 9480 37024
rect 9544 36960 9560 37024
rect 9624 36960 9640 37024
rect 9704 36960 9712 37024
rect 9392 35936 9712 36960
rect 9392 35872 9400 35936
rect 9464 35872 9480 35936
rect 9544 35872 9560 35936
rect 9624 35872 9640 35936
rect 9704 35872 9712 35936
rect 9392 34848 9712 35872
rect 9392 34784 9400 34848
rect 9464 34784 9480 34848
rect 9544 34784 9560 34848
rect 9624 34784 9640 34848
rect 9704 34784 9712 34848
rect 9392 33760 9712 34784
rect 9392 33696 9400 33760
rect 9464 33696 9480 33760
rect 9544 33696 9560 33760
rect 9624 33696 9640 33760
rect 9704 33696 9712 33760
rect 9392 32672 9712 33696
rect 9392 32608 9400 32672
rect 9464 32608 9480 32672
rect 9544 32608 9560 32672
rect 9624 32608 9640 32672
rect 9704 32608 9712 32672
rect 9392 31584 9712 32608
rect 9392 31520 9400 31584
rect 9464 31520 9480 31584
rect 9544 31520 9560 31584
rect 9624 31520 9640 31584
rect 9704 31520 9712 31584
rect 9392 30496 9712 31520
rect 9392 30432 9400 30496
rect 9464 30432 9480 30496
rect 9544 30432 9560 30496
rect 9624 30432 9640 30496
rect 9704 30432 9712 30496
rect 9392 29408 9712 30432
rect 9392 29344 9400 29408
rect 9464 29344 9480 29408
rect 9544 29344 9560 29408
rect 9624 29344 9640 29408
rect 9704 29344 9712 29408
rect 9392 28320 9712 29344
rect 9392 28256 9400 28320
rect 9464 28256 9480 28320
rect 9544 28256 9560 28320
rect 9624 28256 9640 28320
rect 9704 28256 9712 28320
rect 9392 27232 9712 28256
rect 9392 27168 9400 27232
rect 9464 27168 9480 27232
rect 9544 27168 9560 27232
rect 9624 27168 9640 27232
rect 9704 27168 9712 27232
rect 9392 26144 9712 27168
rect 9392 26080 9400 26144
rect 9464 26080 9480 26144
rect 9544 26080 9560 26144
rect 9624 26080 9640 26144
rect 9704 26080 9712 26144
rect 9392 25056 9712 26080
rect 9392 24992 9400 25056
rect 9464 24992 9480 25056
rect 9544 24992 9560 25056
rect 9624 24992 9640 25056
rect 9704 24992 9712 25056
rect 9392 23968 9712 24992
rect 9392 23904 9400 23968
rect 9464 23904 9480 23968
rect 9544 23904 9560 23968
rect 9624 23904 9640 23968
rect 9704 23904 9712 23968
rect 9392 22880 9712 23904
rect 9392 22816 9400 22880
rect 9464 22816 9480 22880
rect 9544 22816 9560 22880
rect 9624 22816 9640 22880
rect 9704 22816 9712 22880
rect 9392 21792 9712 22816
rect 9392 21728 9400 21792
rect 9464 21728 9480 21792
rect 9544 21728 9560 21792
rect 9624 21728 9640 21792
rect 9704 21728 9712 21792
rect 9392 20704 9712 21728
rect 9392 20640 9400 20704
rect 9464 20640 9480 20704
rect 9544 20640 9560 20704
rect 9624 20640 9640 20704
rect 9704 20640 9712 20704
rect 9392 19616 9712 20640
rect 9392 19552 9400 19616
rect 9464 19552 9480 19616
rect 9544 19552 9560 19616
rect 9624 19552 9640 19616
rect 9704 19552 9712 19616
rect 9392 18528 9712 19552
rect 9392 18464 9400 18528
rect 9464 18464 9480 18528
rect 9544 18464 9560 18528
rect 9624 18464 9640 18528
rect 9704 18464 9712 18528
rect 9392 17440 9712 18464
rect 9392 17376 9400 17440
rect 9464 17376 9480 17440
rect 9544 17376 9560 17440
rect 9624 17376 9640 17440
rect 9704 17376 9712 17440
rect 9392 16352 9712 17376
rect 9392 16288 9400 16352
rect 9464 16288 9480 16352
rect 9544 16288 9560 16352
rect 9624 16288 9640 16352
rect 9704 16288 9712 16352
rect 9392 15264 9712 16288
rect 9392 15200 9400 15264
rect 9464 15200 9480 15264
rect 9544 15200 9560 15264
rect 9624 15200 9640 15264
rect 9704 15200 9712 15264
rect 9392 14176 9712 15200
rect 9392 14112 9400 14176
rect 9464 14112 9480 14176
rect 9544 14112 9560 14176
rect 9624 14112 9640 14176
rect 9704 14112 9712 14176
rect 9392 13088 9712 14112
rect 9392 13024 9400 13088
rect 9464 13024 9480 13088
rect 9544 13024 9560 13088
rect 9624 13024 9640 13088
rect 9704 13024 9712 13088
rect 9392 12000 9712 13024
rect 9392 11936 9400 12000
rect 9464 11936 9480 12000
rect 9544 11936 9560 12000
rect 9624 11936 9640 12000
rect 9704 11936 9712 12000
rect 9392 10912 9712 11936
rect 9392 10848 9400 10912
rect 9464 10848 9480 10912
rect 9544 10848 9560 10912
rect 9624 10848 9640 10912
rect 9704 10848 9712 10912
rect 9392 9824 9712 10848
rect 9392 9760 9400 9824
rect 9464 9760 9480 9824
rect 9544 9760 9560 9824
rect 9624 9760 9640 9824
rect 9704 9760 9712 9824
rect 9392 8736 9712 9760
rect 9392 8672 9400 8736
rect 9464 8672 9480 8736
rect 9544 8672 9560 8736
rect 9624 8672 9640 8736
rect 9704 8672 9712 8736
rect 9392 7648 9712 8672
rect 9392 7584 9400 7648
rect 9464 7584 9480 7648
rect 9544 7584 9560 7648
rect 9624 7584 9640 7648
rect 9704 7584 9712 7648
rect 9392 6560 9712 7584
rect 9392 6496 9400 6560
rect 9464 6496 9480 6560
rect 9544 6496 9560 6560
rect 9624 6496 9640 6560
rect 9704 6496 9712 6560
rect 9392 5472 9712 6496
rect 9392 5408 9400 5472
rect 9464 5408 9480 5472
rect 9544 5408 9560 5472
rect 9624 5408 9640 5472
rect 9704 5408 9712 5472
rect 9392 4384 9712 5408
rect 9392 4320 9400 4384
rect 9464 4320 9480 4384
rect 9544 4320 9560 4384
rect 9624 4320 9640 4384
rect 9704 4320 9712 4384
rect 9392 3296 9712 4320
rect 9392 3232 9400 3296
rect 9464 3232 9480 3296
rect 9544 3232 9560 3296
rect 9624 3232 9640 3296
rect 9704 3232 9712 3296
rect 9392 2208 9712 3232
rect 9392 2144 9400 2208
rect 9464 2144 9480 2208
rect 9544 2144 9560 2208
rect 9624 2144 9640 2208
rect 9704 2144 9712 2208
rect 9392 2128 9712 2144
rect 13616 39744 13936 39760
rect 13616 39680 13624 39744
rect 13688 39680 13704 39744
rect 13768 39680 13784 39744
rect 13848 39680 13864 39744
rect 13928 39680 13936 39744
rect 13616 38656 13936 39680
rect 13616 38592 13624 38656
rect 13688 38592 13704 38656
rect 13768 38592 13784 38656
rect 13848 38592 13864 38656
rect 13928 38592 13936 38656
rect 13616 37568 13936 38592
rect 13616 37504 13624 37568
rect 13688 37504 13704 37568
rect 13768 37504 13784 37568
rect 13848 37504 13864 37568
rect 13928 37504 13936 37568
rect 13616 36480 13936 37504
rect 13616 36416 13624 36480
rect 13688 36416 13704 36480
rect 13768 36416 13784 36480
rect 13848 36416 13864 36480
rect 13928 36416 13936 36480
rect 13616 35392 13936 36416
rect 13616 35328 13624 35392
rect 13688 35328 13704 35392
rect 13768 35328 13784 35392
rect 13848 35328 13864 35392
rect 13928 35328 13936 35392
rect 13616 34304 13936 35328
rect 13616 34240 13624 34304
rect 13688 34240 13704 34304
rect 13768 34240 13784 34304
rect 13848 34240 13864 34304
rect 13928 34240 13936 34304
rect 13616 33216 13936 34240
rect 13616 33152 13624 33216
rect 13688 33152 13704 33216
rect 13768 33152 13784 33216
rect 13848 33152 13864 33216
rect 13928 33152 13936 33216
rect 13616 32128 13936 33152
rect 13616 32064 13624 32128
rect 13688 32064 13704 32128
rect 13768 32064 13784 32128
rect 13848 32064 13864 32128
rect 13928 32064 13936 32128
rect 13616 31040 13936 32064
rect 13616 30976 13624 31040
rect 13688 30976 13704 31040
rect 13768 30976 13784 31040
rect 13848 30976 13864 31040
rect 13928 30976 13936 31040
rect 13616 29952 13936 30976
rect 13616 29888 13624 29952
rect 13688 29888 13704 29952
rect 13768 29888 13784 29952
rect 13848 29888 13864 29952
rect 13928 29888 13936 29952
rect 13616 28864 13936 29888
rect 13616 28800 13624 28864
rect 13688 28800 13704 28864
rect 13768 28800 13784 28864
rect 13848 28800 13864 28864
rect 13928 28800 13936 28864
rect 13616 27776 13936 28800
rect 13616 27712 13624 27776
rect 13688 27712 13704 27776
rect 13768 27712 13784 27776
rect 13848 27712 13864 27776
rect 13928 27712 13936 27776
rect 13616 26688 13936 27712
rect 13616 26624 13624 26688
rect 13688 26624 13704 26688
rect 13768 26624 13784 26688
rect 13848 26624 13864 26688
rect 13928 26624 13936 26688
rect 13616 25600 13936 26624
rect 13616 25536 13624 25600
rect 13688 25536 13704 25600
rect 13768 25536 13784 25600
rect 13848 25536 13864 25600
rect 13928 25536 13936 25600
rect 13616 24512 13936 25536
rect 13616 24448 13624 24512
rect 13688 24448 13704 24512
rect 13768 24448 13784 24512
rect 13848 24448 13864 24512
rect 13928 24448 13936 24512
rect 13616 23424 13936 24448
rect 13616 23360 13624 23424
rect 13688 23360 13704 23424
rect 13768 23360 13784 23424
rect 13848 23360 13864 23424
rect 13928 23360 13936 23424
rect 13616 22336 13936 23360
rect 13616 22272 13624 22336
rect 13688 22272 13704 22336
rect 13768 22272 13784 22336
rect 13848 22272 13864 22336
rect 13928 22272 13936 22336
rect 13616 21248 13936 22272
rect 13616 21184 13624 21248
rect 13688 21184 13704 21248
rect 13768 21184 13784 21248
rect 13848 21184 13864 21248
rect 13928 21184 13936 21248
rect 13616 20160 13936 21184
rect 13616 20096 13624 20160
rect 13688 20096 13704 20160
rect 13768 20096 13784 20160
rect 13848 20096 13864 20160
rect 13928 20096 13936 20160
rect 13616 19072 13936 20096
rect 13616 19008 13624 19072
rect 13688 19008 13704 19072
rect 13768 19008 13784 19072
rect 13848 19008 13864 19072
rect 13928 19008 13936 19072
rect 13616 17984 13936 19008
rect 13616 17920 13624 17984
rect 13688 17920 13704 17984
rect 13768 17920 13784 17984
rect 13848 17920 13864 17984
rect 13928 17920 13936 17984
rect 13616 16896 13936 17920
rect 13616 16832 13624 16896
rect 13688 16832 13704 16896
rect 13768 16832 13784 16896
rect 13848 16832 13864 16896
rect 13928 16832 13936 16896
rect 13616 15808 13936 16832
rect 13616 15744 13624 15808
rect 13688 15744 13704 15808
rect 13768 15744 13784 15808
rect 13848 15744 13864 15808
rect 13928 15744 13936 15808
rect 13616 14720 13936 15744
rect 13616 14656 13624 14720
rect 13688 14656 13704 14720
rect 13768 14656 13784 14720
rect 13848 14656 13864 14720
rect 13928 14656 13936 14720
rect 13616 13632 13936 14656
rect 13616 13568 13624 13632
rect 13688 13568 13704 13632
rect 13768 13568 13784 13632
rect 13848 13568 13864 13632
rect 13928 13568 13936 13632
rect 13616 12544 13936 13568
rect 13616 12480 13624 12544
rect 13688 12480 13704 12544
rect 13768 12480 13784 12544
rect 13848 12480 13864 12544
rect 13928 12480 13936 12544
rect 13616 11456 13936 12480
rect 13616 11392 13624 11456
rect 13688 11392 13704 11456
rect 13768 11392 13784 11456
rect 13848 11392 13864 11456
rect 13928 11392 13936 11456
rect 13616 10368 13936 11392
rect 13616 10304 13624 10368
rect 13688 10304 13704 10368
rect 13768 10304 13784 10368
rect 13848 10304 13864 10368
rect 13928 10304 13936 10368
rect 13616 9280 13936 10304
rect 13616 9216 13624 9280
rect 13688 9216 13704 9280
rect 13768 9216 13784 9280
rect 13848 9216 13864 9280
rect 13928 9216 13936 9280
rect 13616 8192 13936 9216
rect 13616 8128 13624 8192
rect 13688 8128 13704 8192
rect 13768 8128 13784 8192
rect 13848 8128 13864 8192
rect 13928 8128 13936 8192
rect 13616 7104 13936 8128
rect 13616 7040 13624 7104
rect 13688 7040 13704 7104
rect 13768 7040 13784 7104
rect 13848 7040 13864 7104
rect 13928 7040 13936 7104
rect 13616 6016 13936 7040
rect 13616 5952 13624 6016
rect 13688 5952 13704 6016
rect 13768 5952 13784 6016
rect 13848 5952 13864 6016
rect 13928 5952 13936 6016
rect 13616 4928 13936 5952
rect 13616 4864 13624 4928
rect 13688 4864 13704 4928
rect 13768 4864 13784 4928
rect 13848 4864 13864 4928
rect 13928 4864 13936 4928
rect 13616 3840 13936 4864
rect 13616 3776 13624 3840
rect 13688 3776 13704 3840
rect 13768 3776 13784 3840
rect 13848 3776 13864 3840
rect 13928 3776 13936 3840
rect 13616 2752 13936 3776
rect 13616 2688 13624 2752
rect 13688 2688 13704 2752
rect 13768 2688 13784 2752
rect 13848 2688 13864 2752
rect 13928 2688 13936 2752
rect 13616 2128 13936 2688
rect 17840 39200 18160 39760
rect 17840 39136 17848 39200
rect 17912 39136 17928 39200
rect 17992 39136 18008 39200
rect 18072 39136 18088 39200
rect 18152 39136 18160 39200
rect 17840 38112 18160 39136
rect 17840 38048 17848 38112
rect 17912 38048 17928 38112
rect 17992 38048 18008 38112
rect 18072 38048 18088 38112
rect 18152 38048 18160 38112
rect 17840 37024 18160 38048
rect 17840 36960 17848 37024
rect 17912 36960 17928 37024
rect 17992 36960 18008 37024
rect 18072 36960 18088 37024
rect 18152 36960 18160 37024
rect 17840 35936 18160 36960
rect 17840 35872 17848 35936
rect 17912 35872 17928 35936
rect 17992 35872 18008 35936
rect 18072 35872 18088 35936
rect 18152 35872 18160 35936
rect 17840 34848 18160 35872
rect 17840 34784 17848 34848
rect 17912 34784 17928 34848
rect 17992 34784 18008 34848
rect 18072 34784 18088 34848
rect 18152 34784 18160 34848
rect 17840 33760 18160 34784
rect 17840 33696 17848 33760
rect 17912 33696 17928 33760
rect 17992 33696 18008 33760
rect 18072 33696 18088 33760
rect 18152 33696 18160 33760
rect 17840 32672 18160 33696
rect 17840 32608 17848 32672
rect 17912 32608 17928 32672
rect 17992 32608 18008 32672
rect 18072 32608 18088 32672
rect 18152 32608 18160 32672
rect 17840 31584 18160 32608
rect 17840 31520 17848 31584
rect 17912 31520 17928 31584
rect 17992 31520 18008 31584
rect 18072 31520 18088 31584
rect 18152 31520 18160 31584
rect 17840 30496 18160 31520
rect 17840 30432 17848 30496
rect 17912 30432 17928 30496
rect 17992 30432 18008 30496
rect 18072 30432 18088 30496
rect 18152 30432 18160 30496
rect 17840 29408 18160 30432
rect 17840 29344 17848 29408
rect 17912 29344 17928 29408
rect 17992 29344 18008 29408
rect 18072 29344 18088 29408
rect 18152 29344 18160 29408
rect 17840 28320 18160 29344
rect 17840 28256 17848 28320
rect 17912 28256 17928 28320
rect 17992 28256 18008 28320
rect 18072 28256 18088 28320
rect 18152 28256 18160 28320
rect 17840 27232 18160 28256
rect 17840 27168 17848 27232
rect 17912 27168 17928 27232
rect 17992 27168 18008 27232
rect 18072 27168 18088 27232
rect 18152 27168 18160 27232
rect 17840 26144 18160 27168
rect 17840 26080 17848 26144
rect 17912 26080 17928 26144
rect 17992 26080 18008 26144
rect 18072 26080 18088 26144
rect 18152 26080 18160 26144
rect 17840 25056 18160 26080
rect 17840 24992 17848 25056
rect 17912 24992 17928 25056
rect 17992 24992 18008 25056
rect 18072 24992 18088 25056
rect 18152 24992 18160 25056
rect 17840 23968 18160 24992
rect 17840 23904 17848 23968
rect 17912 23904 17928 23968
rect 17992 23904 18008 23968
rect 18072 23904 18088 23968
rect 18152 23904 18160 23968
rect 17840 22880 18160 23904
rect 17840 22816 17848 22880
rect 17912 22816 17928 22880
rect 17992 22816 18008 22880
rect 18072 22816 18088 22880
rect 18152 22816 18160 22880
rect 17840 21792 18160 22816
rect 17840 21728 17848 21792
rect 17912 21728 17928 21792
rect 17992 21728 18008 21792
rect 18072 21728 18088 21792
rect 18152 21728 18160 21792
rect 17840 20704 18160 21728
rect 17840 20640 17848 20704
rect 17912 20640 17928 20704
rect 17992 20640 18008 20704
rect 18072 20640 18088 20704
rect 18152 20640 18160 20704
rect 17840 19616 18160 20640
rect 17840 19552 17848 19616
rect 17912 19552 17928 19616
rect 17992 19552 18008 19616
rect 18072 19552 18088 19616
rect 18152 19552 18160 19616
rect 17840 18528 18160 19552
rect 17840 18464 17848 18528
rect 17912 18464 17928 18528
rect 17992 18464 18008 18528
rect 18072 18464 18088 18528
rect 18152 18464 18160 18528
rect 17840 17440 18160 18464
rect 17840 17376 17848 17440
rect 17912 17376 17928 17440
rect 17992 17376 18008 17440
rect 18072 17376 18088 17440
rect 18152 17376 18160 17440
rect 17840 16352 18160 17376
rect 17840 16288 17848 16352
rect 17912 16288 17928 16352
rect 17992 16288 18008 16352
rect 18072 16288 18088 16352
rect 18152 16288 18160 16352
rect 17840 15264 18160 16288
rect 17840 15200 17848 15264
rect 17912 15200 17928 15264
rect 17992 15200 18008 15264
rect 18072 15200 18088 15264
rect 18152 15200 18160 15264
rect 17840 14176 18160 15200
rect 17840 14112 17848 14176
rect 17912 14112 17928 14176
rect 17992 14112 18008 14176
rect 18072 14112 18088 14176
rect 18152 14112 18160 14176
rect 17840 13088 18160 14112
rect 17840 13024 17848 13088
rect 17912 13024 17928 13088
rect 17992 13024 18008 13088
rect 18072 13024 18088 13088
rect 18152 13024 18160 13088
rect 17840 12000 18160 13024
rect 17840 11936 17848 12000
rect 17912 11936 17928 12000
rect 17992 11936 18008 12000
rect 18072 11936 18088 12000
rect 18152 11936 18160 12000
rect 17840 10912 18160 11936
rect 17840 10848 17848 10912
rect 17912 10848 17928 10912
rect 17992 10848 18008 10912
rect 18072 10848 18088 10912
rect 18152 10848 18160 10912
rect 17840 9824 18160 10848
rect 17840 9760 17848 9824
rect 17912 9760 17928 9824
rect 17992 9760 18008 9824
rect 18072 9760 18088 9824
rect 18152 9760 18160 9824
rect 17840 8736 18160 9760
rect 17840 8672 17848 8736
rect 17912 8672 17928 8736
rect 17992 8672 18008 8736
rect 18072 8672 18088 8736
rect 18152 8672 18160 8736
rect 17840 7648 18160 8672
rect 17840 7584 17848 7648
rect 17912 7584 17928 7648
rect 17992 7584 18008 7648
rect 18072 7584 18088 7648
rect 18152 7584 18160 7648
rect 17840 6560 18160 7584
rect 17840 6496 17848 6560
rect 17912 6496 17928 6560
rect 17992 6496 18008 6560
rect 18072 6496 18088 6560
rect 18152 6496 18160 6560
rect 17840 5472 18160 6496
rect 17840 5408 17848 5472
rect 17912 5408 17928 5472
rect 17992 5408 18008 5472
rect 18072 5408 18088 5472
rect 18152 5408 18160 5472
rect 17840 4384 18160 5408
rect 17840 4320 17848 4384
rect 17912 4320 17928 4384
rect 17992 4320 18008 4384
rect 18072 4320 18088 4384
rect 18152 4320 18160 4384
rect 17840 3296 18160 4320
rect 17840 3232 17848 3296
rect 17912 3232 17928 3296
rect 17992 3232 18008 3296
rect 18072 3232 18088 3296
rect 18152 3232 18160 3296
rect 17840 2208 18160 3232
rect 17840 2144 17848 2208
rect 17912 2144 17928 2208
rect 17992 2144 18008 2208
rect 18072 2144 18088 2208
rect 18152 2144 18160 2208
rect 17840 2128 18160 2144
rect 22064 39744 22384 39760
rect 22064 39680 22072 39744
rect 22136 39680 22152 39744
rect 22216 39680 22232 39744
rect 22296 39680 22312 39744
rect 22376 39680 22384 39744
rect 22064 38656 22384 39680
rect 22064 38592 22072 38656
rect 22136 38592 22152 38656
rect 22216 38592 22232 38656
rect 22296 38592 22312 38656
rect 22376 38592 22384 38656
rect 22064 37568 22384 38592
rect 22064 37504 22072 37568
rect 22136 37504 22152 37568
rect 22216 37504 22232 37568
rect 22296 37504 22312 37568
rect 22376 37504 22384 37568
rect 22064 36480 22384 37504
rect 22064 36416 22072 36480
rect 22136 36416 22152 36480
rect 22216 36416 22232 36480
rect 22296 36416 22312 36480
rect 22376 36416 22384 36480
rect 22064 35392 22384 36416
rect 22064 35328 22072 35392
rect 22136 35328 22152 35392
rect 22216 35328 22232 35392
rect 22296 35328 22312 35392
rect 22376 35328 22384 35392
rect 22064 34304 22384 35328
rect 22064 34240 22072 34304
rect 22136 34240 22152 34304
rect 22216 34240 22232 34304
rect 22296 34240 22312 34304
rect 22376 34240 22384 34304
rect 22064 33216 22384 34240
rect 22064 33152 22072 33216
rect 22136 33152 22152 33216
rect 22216 33152 22232 33216
rect 22296 33152 22312 33216
rect 22376 33152 22384 33216
rect 22064 32128 22384 33152
rect 22064 32064 22072 32128
rect 22136 32064 22152 32128
rect 22216 32064 22232 32128
rect 22296 32064 22312 32128
rect 22376 32064 22384 32128
rect 22064 31040 22384 32064
rect 22064 30976 22072 31040
rect 22136 30976 22152 31040
rect 22216 30976 22232 31040
rect 22296 30976 22312 31040
rect 22376 30976 22384 31040
rect 22064 29952 22384 30976
rect 22064 29888 22072 29952
rect 22136 29888 22152 29952
rect 22216 29888 22232 29952
rect 22296 29888 22312 29952
rect 22376 29888 22384 29952
rect 22064 28864 22384 29888
rect 22064 28800 22072 28864
rect 22136 28800 22152 28864
rect 22216 28800 22232 28864
rect 22296 28800 22312 28864
rect 22376 28800 22384 28864
rect 22064 27776 22384 28800
rect 22064 27712 22072 27776
rect 22136 27712 22152 27776
rect 22216 27712 22232 27776
rect 22296 27712 22312 27776
rect 22376 27712 22384 27776
rect 22064 26688 22384 27712
rect 22064 26624 22072 26688
rect 22136 26624 22152 26688
rect 22216 26624 22232 26688
rect 22296 26624 22312 26688
rect 22376 26624 22384 26688
rect 22064 25600 22384 26624
rect 22064 25536 22072 25600
rect 22136 25536 22152 25600
rect 22216 25536 22232 25600
rect 22296 25536 22312 25600
rect 22376 25536 22384 25600
rect 22064 24512 22384 25536
rect 22064 24448 22072 24512
rect 22136 24448 22152 24512
rect 22216 24448 22232 24512
rect 22296 24448 22312 24512
rect 22376 24448 22384 24512
rect 22064 23424 22384 24448
rect 22064 23360 22072 23424
rect 22136 23360 22152 23424
rect 22216 23360 22232 23424
rect 22296 23360 22312 23424
rect 22376 23360 22384 23424
rect 22064 22336 22384 23360
rect 22064 22272 22072 22336
rect 22136 22272 22152 22336
rect 22216 22272 22232 22336
rect 22296 22272 22312 22336
rect 22376 22272 22384 22336
rect 22064 21248 22384 22272
rect 22064 21184 22072 21248
rect 22136 21184 22152 21248
rect 22216 21184 22232 21248
rect 22296 21184 22312 21248
rect 22376 21184 22384 21248
rect 22064 20160 22384 21184
rect 22064 20096 22072 20160
rect 22136 20096 22152 20160
rect 22216 20096 22232 20160
rect 22296 20096 22312 20160
rect 22376 20096 22384 20160
rect 22064 19072 22384 20096
rect 22064 19008 22072 19072
rect 22136 19008 22152 19072
rect 22216 19008 22232 19072
rect 22296 19008 22312 19072
rect 22376 19008 22384 19072
rect 22064 17984 22384 19008
rect 22064 17920 22072 17984
rect 22136 17920 22152 17984
rect 22216 17920 22232 17984
rect 22296 17920 22312 17984
rect 22376 17920 22384 17984
rect 22064 16896 22384 17920
rect 22064 16832 22072 16896
rect 22136 16832 22152 16896
rect 22216 16832 22232 16896
rect 22296 16832 22312 16896
rect 22376 16832 22384 16896
rect 22064 15808 22384 16832
rect 22064 15744 22072 15808
rect 22136 15744 22152 15808
rect 22216 15744 22232 15808
rect 22296 15744 22312 15808
rect 22376 15744 22384 15808
rect 22064 14720 22384 15744
rect 22064 14656 22072 14720
rect 22136 14656 22152 14720
rect 22216 14656 22232 14720
rect 22296 14656 22312 14720
rect 22376 14656 22384 14720
rect 22064 13632 22384 14656
rect 22064 13568 22072 13632
rect 22136 13568 22152 13632
rect 22216 13568 22232 13632
rect 22296 13568 22312 13632
rect 22376 13568 22384 13632
rect 22064 12544 22384 13568
rect 22064 12480 22072 12544
rect 22136 12480 22152 12544
rect 22216 12480 22232 12544
rect 22296 12480 22312 12544
rect 22376 12480 22384 12544
rect 22064 11456 22384 12480
rect 22064 11392 22072 11456
rect 22136 11392 22152 11456
rect 22216 11392 22232 11456
rect 22296 11392 22312 11456
rect 22376 11392 22384 11456
rect 22064 10368 22384 11392
rect 22064 10304 22072 10368
rect 22136 10304 22152 10368
rect 22216 10304 22232 10368
rect 22296 10304 22312 10368
rect 22376 10304 22384 10368
rect 22064 9280 22384 10304
rect 22064 9216 22072 9280
rect 22136 9216 22152 9280
rect 22216 9216 22232 9280
rect 22296 9216 22312 9280
rect 22376 9216 22384 9280
rect 22064 8192 22384 9216
rect 22064 8128 22072 8192
rect 22136 8128 22152 8192
rect 22216 8128 22232 8192
rect 22296 8128 22312 8192
rect 22376 8128 22384 8192
rect 22064 7104 22384 8128
rect 22064 7040 22072 7104
rect 22136 7040 22152 7104
rect 22216 7040 22232 7104
rect 22296 7040 22312 7104
rect 22376 7040 22384 7104
rect 22064 6016 22384 7040
rect 22064 5952 22072 6016
rect 22136 5952 22152 6016
rect 22216 5952 22232 6016
rect 22296 5952 22312 6016
rect 22376 5952 22384 6016
rect 22064 4928 22384 5952
rect 22064 4864 22072 4928
rect 22136 4864 22152 4928
rect 22216 4864 22232 4928
rect 22296 4864 22312 4928
rect 22376 4864 22384 4928
rect 22064 3840 22384 4864
rect 22064 3776 22072 3840
rect 22136 3776 22152 3840
rect 22216 3776 22232 3840
rect 22296 3776 22312 3840
rect 22376 3776 22384 3840
rect 22064 2752 22384 3776
rect 22064 2688 22072 2752
rect 22136 2688 22152 2752
rect 22216 2688 22232 2752
rect 22296 2688 22312 2752
rect 22376 2688 22384 2752
rect 22064 2128 22384 2688
rect 26288 39200 26608 39760
rect 26288 39136 26296 39200
rect 26360 39136 26376 39200
rect 26440 39136 26456 39200
rect 26520 39136 26536 39200
rect 26600 39136 26608 39200
rect 26288 38112 26608 39136
rect 26288 38048 26296 38112
rect 26360 38048 26376 38112
rect 26440 38048 26456 38112
rect 26520 38048 26536 38112
rect 26600 38048 26608 38112
rect 26288 37024 26608 38048
rect 26288 36960 26296 37024
rect 26360 36960 26376 37024
rect 26440 36960 26456 37024
rect 26520 36960 26536 37024
rect 26600 36960 26608 37024
rect 26288 35936 26608 36960
rect 26288 35872 26296 35936
rect 26360 35872 26376 35936
rect 26440 35872 26456 35936
rect 26520 35872 26536 35936
rect 26600 35872 26608 35936
rect 26288 34848 26608 35872
rect 26288 34784 26296 34848
rect 26360 34784 26376 34848
rect 26440 34784 26456 34848
rect 26520 34784 26536 34848
rect 26600 34784 26608 34848
rect 26288 33760 26608 34784
rect 26288 33696 26296 33760
rect 26360 33696 26376 33760
rect 26440 33696 26456 33760
rect 26520 33696 26536 33760
rect 26600 33696 26608 33760
rect 26288 32672 26608 33696
rect 26288 32608 26296 32672
rect 26360 32608 26376 32672
rect 26440 32608 26456 32672
rect 26520 32608 26536 32672
rect 26600 32608 26608 32672
rect 26288 31584 26608 32608
rect 26288 31520 26296 31584
rect 26360 31520 26376 31584
rect 26440 31520 26456 31584
rect 26520 31520 26536 31584
rect 26600 31520 26608 31584
rect 26288 30496 26608 31520
rect 26288 30432 26296 30496
rect 26360 30432 26376 30496
rect 26440 30432 26456 30496
rect 26520 30432 26536 30496
rect 26600 30432 26608 30496
rect 26288 29408 26608 30432
rect 26288 29344 26296 29408
rect 26360 29344 26376 29408
rect 26440 29344 26456 29408
rect 26520 29344 26536 29408
rect 26600 29344 26608 29408
rect 26288 28320 26608 29344
rect 26288 28256 26296 28320
rect 26360 28256 26376 28320
rect 26440 28256 26456 28320
rect 26520 28256 26536 28320
rect 26600 28256 26608 28320
rect 26288 27232 26608 28256
rect 26288 27168 26296 27232
rect 26360 27168 26376 27232
rect 26440 27168 26456 27232
rect 26520 27168 26536 27232
rect 26600 27168 26608 27232
rect 26288 26144 26608 27168
rect 26288 26080 26296 26144
rect 26360 26080 26376 26144
rect 26440 26080 26456 26144
rect 26520 26080 26536 26144
rect 26600 26080 26608 26144
rect 26288 25056 26608 26080
rect 26288 24992 26296 25056
rect 26360 24992 26376 25056
rect 26440 24992 26456 25056
rect 26520 24992 26536 25056
rect 26600 24992 26608 25056
rect 26288 23968 26608 24992
rect 26288 23904 26296 23968
rect 26360 23904 26376 23968
rect 26440 23904 26456 23968
rect 26520 23904 26536 23968
rect 26600 23904 26608 23968
rect 26288 22880 26608 23904
rect 26288 22816 26296 22880
rect 26360 22816 26376 22880
rect 26440 22816 26456 22880
rect 26520 22816 26536 22880
rect 26600 22816 26608 22880
rect 26288 21792 26608 22816
rect 26288 21728 26296 21792
rect 26360 21728 26376 21792
rect 26440 21728 26456 21792
rect 26520 21728 26536 21792
rect 26600 21728 26608 21792
rect 26288 20704 26608 21728
rect 26288 20640 26296 20704
rect 26360 20640 26376 20704
rect 26440 20640 26456 20704
rect 26520 20640 26536 20704
rect 26600 20640 26608 20704
rect 26288 19616 26608 20640
rect 26288 19552 26296 19616
rect 26360 19552 26376 19616
rect 26440 19552 26456 19616
rect 26520 19552 26536 19616
rect 26600 19552 26608 19616
rect 26288 18528 26608 19552
rect 26288 18464 26296 18528
rect 26360 18464 26376 18528
rect 26440 18464 26456 18528
rect 26520 18464 26536 18528
rect 26600 18464 26608 18528
rect 26288 17440 26608 18464
rect 26288 17376 26296 17440
rect 26360 17376 26376 17440
rect 26440 17376 26456 17440
rect 26520 17376 26536 17440
rect 26600 17376 26608 17440
rect 26288 16352 26608 17376
rect 26288 16288 26296 16352
rect 26360 16288 26376 16352
rect 26440 16288 26456 16352
rect 26520 16288 26536 16352
rect 26600 16288 26608 16352
rect 26288 15264 26608 16288
rect 26288 15200 26296 15264
rect 26360 15200 26376 15264
rect 26440 15200 26456 15264
rect 26520 15200 26536 15264
rect 26600 15200 26608 15264
rect 26288 14176 26608 15200
rect 26288 14112 26296 14176
rect 26360 14112 26376 14176
rect 26440 14112 26456 14176
rect 26520 14112 26536 14176
rect 26600 14112 26608 14176
rect 26288 13088 26608 14112
rect 26288 13024 26296 13088
rect 26360 13024 26376 13088
rect 26440 13024 26456 13088
rect 26520 13024 26536 13088
rect 26600 13024 26608 13088
rect 26288 12000 26608 13024
rect 26288 11936 26296 12000
rect 26360 11936 26376 12000
rect 26440 11936 26456 12000
rect 26520 11936 26536 12000
rect 26600 11936 26608 12000
rect 26288 10912 26608 11936
rect 26288 10848 26296 10912
rect 26360 10848 26376 10912
rect 26440 10848 26456 10912
rect 26520 10848 26536 10912
rect 26600 10848 26608 10912
rect 26288 9824 26608 10848
rect 26288 9760 26296 9824
rect 26360 9760 26376 9824
rect 26440 9760 26456 9824
rect 26520 9760 26536 9824
rect 26600 9760 26608 9824
rect 26288 8736 26608 9760
rect 26288 8672 26296 8736
rect 26360 8672 26376 8736
rect 26440 8672 26456 8736
rect 26520 8672 26536 8736
rect 26600 8672 26608 8736
rect 26288 7648 26608 8672
rect 26288 7584 26296 7648
rect 26360 7584 26376 7648
rect 26440 7584 26456 7648
rect 26520 7584 26536 7648
rect 26600 7584 26608 7648
rect 26288 6560 26608 7584
rect 26288 6496 26296 6560
rect 26360 6496 26376 6560
rect 26440 6496 26456 6560
rect 26520 6496 26536 6560
rect 26600 6496 26608 6560
rect 26288 5472 26608 6496
rect 26288 5408 26296 5472
rect 26360 5408 26376 5472
rect 26440 5408 26456 5472
rect 26520 5408 26536 5472
rect 26600 5408 26608 5472
rect 26288 4384 26608 5408
rect 26288 4320 26296 4384
rect 26360 4320 26376 4384
rect 26440 4320 26456 4384
rect 26520 4320 26536 4384
rect 26600 4320 26608 4384
rect 26288 3296 26608 4320
rect 26288 3232 26296 3296
rect 26360 3232 26376 3296
rect 26440 3232 26456 3296
rect 26520 3232 26536 3296
rect 26600 3232 26608 3296
rect 26288 2208 26608 3232
rect 26288 2144 26296 2208
rect 26360 2144 26376 2208
rect 26440 2144 26456 2208
rect 26520 2144 26536 2208
rect 26600 2144 26608 2208
rect 26288 2128 26608 2144
rect 30512 39744 30832 39760
rect 30512 39680 30520 39744
rect 30584 39680 30600 39744
rect 30664 39680 30680 39744
rect 30744 39680 30760 39744
rect 30824 39680 30832 39744
rect 30512 38656 30832 39680
rect 30512 38592 30520 38656
rect 30584 38592 30600 38656
rect 30664 38592 30680 38656
rect 30744 38592 30760 38656
rect 30824 38592 30832 38656
rect 30512 37568 30832 38592
rect 30512 37504 30520 37568
rect 30584 37504 30600 37568
rect 30664 37504 30680 37568
rect 30744 37504 30760 37568
rect 30824 37504 30832 37568
rect 30512 36480 30832 37504
rect 30512 36416 30520 36480
rect 30584 36416 30600 36480
rect 30664 36416 30680 36480
rect 30744 36416 30760 36480
rect 30824 36416 30832 36480
rect 30512 35392 30832 36416
rect 30512 35328 30520 35392
rect 30584 35328 30600 35392
rect 30664 35328 30680 35392
rect 30744 35328 30760 35392
rect 30824 35328 30832 35392
rect 30512 34304 30832 35328
rect 30512 34240 30520 34304
rect 30584 34240 30600 34304
rect 30664 34240 30680 34304
rect 30744 34240 30760 34304
rect 30824 34240 30832 34304
rect 30512 33216 30832 34240
rect 30512 33152 30520 33216
rect 30584 33152 30600 33216
rect 30664 33152 30680 33216
rect 30744 33152 30760 33216
rect 30824 33152 30832 33216
rect 30512 32128 30832 33152
rect 30512 32064 30520 32128
rect 30584 32064 30600 32128
rect 30664 32064 30680 32128
rect 30744 32064 30760 32128
rect 30824 32064 30832 32128
rect 30512 31040 30832 32064
rect 30512 30976 30520 31040
rect 30584 30976 30600 31040
rect 30664 30976 30680 31040
rect 30744 30976 30760 31040
rect 30824 30976 30832 31040
rect 30512 29952 30832 30976
rect 30512 29888 30520 29952
rect 30584 29888 30600 29952
rect 30664 29888 30680 29952
rect 30744 29888 30760 29952
rect 30824 29888 30832 29952
rect 30512 28864 30832 29888
rect 30512 28800 30520 28864
rect 30584 28800 30600 28864
rect 30664 28800 30680 28864
rect 30744 28800 30760 28864
rect 30824 28800 30832 28864
rect 30512 27776 30832 28800
rect 30512 27712 30520 27776
rect 30584 27712 30600 27776
rect 30664 27712 30680 27776
rect 30744 27712 30760 27776
rect 30824 27712 30832 27776
rect 30512 26688 30832 27712
rect 30512 26624 30520 26688
rect 30584 26624 30600 26688
rect 30664 26624 30680 26688
rect 30744 26624 30760 26688
rect 30824 26624 30832 26688
rect 30512 25600 30832 26624
rect 30512 25536 30520 25600
rect 30584 25536 30600 25600
rect 30664 25536 30680 25600
rect 30744 25536 30760 25600
rect 30824 25536 30832 25600
rect 30512 24512 30832 25536
rect 30512 24448 30520 24512
rect 30584 24448 30600 24512
rect 30664 24448 30680 24512
rect 30744 24448 30760 24512
rect 30824 24448 30832 24512
rect 30512 23424 30832 24448
rect 30512 23360 30520 23424
rect 30584 23360 30600 23424
rect 30664 23360 30680 23424
rect 30744 23360 30760 23424
rect 30824 23360 30832 23424
rect 30512 22336 30832 23360
rect 30512 22272 30520 22336
rect 30584 22272 30600 22336
rect 30664 22272 30680 22336
rect 30744 22272 30760 22336
rect 30824 22272 30832 22336
rect 30512 21248 30832 22272
rect 30512 21184 30520 21248
rect 30584 21184 30600 21248
rect 30664 21184 30680 21248
rect 30744 21184 30760 21248
rect 30824 21184 30832 21248
rect 30512 20160 30832 21184
rect 30512 20096 30520 20160
rect 30584 20096 30600 20160
rect 30664 20096 30680 20160
rect 30744 20096 30760 20160
rect 30824 20096 30832 20160
rect 30512 19072 30832 20096
rect 30512 19008 30520 19072
rect 30584 19008 30600 19072
rect 30664 19008 30680 19072
rect 30744 19008 30760 19072
rect 30824 19008 30832 19072
rect 30512 17984 30832 19008
rect 30512 17920 30520 17984
rect 30584 17920 30600 17984
rect 30664 17920 30680 17984
rect 30744 17920 30760 17984
rect 30824 17920 30832 17984
rect 30512 16896 30832 17920
rect 30512 16832 30520 16896
rect 30584 16832 30600 16896
rect 30664 16832 30680 16896
rect 30744 16832 30760 16896
rect 30824 16832 30832 16896
rect 30512 15808 30832 16832
rect 30512 15744 30520 15808
rect 30584 15744 30600 15808
rect 30664 15744 30680 15808
rect 30744 15744 30760 15808
rect 30824 15744 30832 15808
rect 30512 14720 30832 15744
rect 30512 14656 30520 14720
rect 30584 14656 30600 14720
rect 30664 14656 30680 14720
rect 30744 14656 30760 14720
rect 30824 14656 30832 14720
rect 30512 13632 30832 14656
rect 30512 13568 30520 13632
rect 30584 13568 30600 13632
rect 30664 13568 30680 13632
rect 30744 13568 30760 13632
rect 30824 13568 30832 13632
rect 30512 12544 30832 13568
rect 30512 12480 30520 12544
rect 30584 12480 30600 12544
rect 30664 12480 30680 12544
rect 30744 12480 30760 12544
rect 30824 12480 30832 12544
rect 30512 11456 30832 12480
rect 30512 11392 30520 11456
rect 30584 11392 30600 11456
rect 30664 11392 30680 11456
rect 30744 11392 30760 11456
rect 30824 11392 30832 11456
rect 30512 10368 30832 11392
rect 30512 10304 30520 10368
rect 30584 10304 30600 10368
rect 30664 10304 30680 10368
rect 30744 10304 30760 10368
rect 30824 10304 30832 10368
rect 30512 9280 30832 10304
rect 30512 9216 30520 9280
rect 30584 9216 30600 9280
rect 30664 9216 30680 9280
rect 30744 9216 30760 9280
rect 30824 9216 30832 9280
rect 30512 8192 30832 9216
rect 30512 8128 30520 8192
rect 30584 8128 30600 8192
rect 30664 8128 30680 8192
rect 30744 8128 30760 8192
rect 30824 8128 30832 8192
rect 30512 7104 30832 8128
rect 30512 7040 30520 7104
rect 30584 7040 30600 7104
rect 30664 7040 30680 7104
rect 30744 7040 30760 7104
rect 30824 7040 30832 7104
rect 30512 6016 30832 7040
rect 30512 5952 30520 6016
rect 30584 5952 30600 6016
rect 30664 5952 30680 6016
rect 30744 5952 30760 6016
rect 30824 5952 30832 6016
rect 30512 4928 30832 5952
rect 30512 4864 30520 4928
rect 30584 4864 30600 4928
rect 30664 4864 30680 4928
rect 30744 4864 30760 4928
rect 30824 4864 30832 4928
rect 30512 3840 30832 4864
rect 30512 3776 30520 3840
rect 30584 3776 30600 3840
rect 30664 3776 30680 3840
rect 30744 3776 30760 3840
rect 30824 3776 30832 3840
rect 30512 2752 30832 3776
rect 30512 2688 30520 2752
rect 30584 2688 30600 2752
rect 30664 2688 30680 2752
rect 30744 2688 30760 2752
rect 30824 2688 30832 2752
rect 30512 2128 30832 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_200
timestamp 1649977179
transform 1 0 19504 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1649977179
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_115
timestamp 1649977179
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_127
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_86
timestamp 1649977179
transform 1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_320
timestamp 1649977179
transform 1 0 30544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1649977179
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_341
timestamp 1649977179
transform 1 0 32476 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_348
timestamp 1649977179
transform 1 0 33120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1649977179
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1649977179
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_283
timestamp 1649977179
transform 1 0 27140 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_287
timestamp 1649977179
transform 1 0 27508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_299
timestamp 1649977179
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_338
timestamp 1649977179
transform 1 0 32200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_350
timestamp 1649977179
transform 1 0 33304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_61
timestamp 1649977179
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_75
timestamp 1649977179
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_116
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_152
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_308
timestamp 1649977179
transform 1 0 29440 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_316
timestamp 1649977179
transform 1 0 30176 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1649977179
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1649977179
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_90
timestamp 1649977179
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_119
timestamp 1649977179
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_162
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_174
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_283
timestamp 1649977179
transform 1 0 27140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_287
timestamp 1649977179
transform 1 0 27508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_291
timestamp 1649977179
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1649977179
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_342
timestamp 1649977179
transform 1 0 32568 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1649977179
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1649977179
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_344
timestamp 1649977179
transform 1 0 32752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_356
timestamp 1649977179
transform 1 0 33856 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1649977179
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1649977179
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_114
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_144
timestamp 1649977179
transform 1 0 14352 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_168
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1649977179
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1649977179
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_283
timestamp 1649977179
transform 1 0 27140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_287
timestamp 1649977179
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1649977179
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_317
timestamp 1649977179
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_323
timestamp 1649977179
transform 1 0 30820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_330
timestamp 1649977179
transform 1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_338
timestamp 1649977179
transform 1 0 32200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_68
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_92
timestamp 1649977179
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1649977179
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1649977179
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_17
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_330
timestamp 1649977179
transform 1 0 31464 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_342
timestamp 1649977179
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_354
timestamp 1649977179
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1649977179
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_123
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_135
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_147
timestamp 1649977179
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1649977179
transform 1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1649977179
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1649977179
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_301
timestamp 1649977179
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1649977179
transform 1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_314
timestamp 1649977179
transform 1 0 29992 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1649977179
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_227
timestamp 1649977179
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_239
timestamp 1649977179
transform 1 0 23092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_256
timestamp 1649977179
transform 1 0 24656 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_268
timestamp 1649977179
transform 1 0 25760 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_280
timestamp 1649977179
transform 1 0 26864 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_292
timestamp 1649977179
transform 1 0 27968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_138
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_150
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1649977179
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1649977179
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_96
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_108
timestamp 1649977179
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_215
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_227
timestamp 1649977179
transform 1 0 21988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_239
timestamp 1649977179
transform 1 0 23092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_294
timestamp 1649977179
transform 1 0 28152 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1649977179
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_11
timestamp 1649977179
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_47
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_60
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_72
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1649977179
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1649977179
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_311
timestamp 1649977179
transform 1 0 29716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_323
timestamp 1649977179
transform 1 0 30820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_68
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_91
timestamp 1649977179
transform 1 0 9476 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_103
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_115
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_234
timestamp 1649977179
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1649977179
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_146
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_180
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_192
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1649977179
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_344
timestamp 1649977179
transform 1 0 32752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_352
timestamp 1649977179
transform 1 0 33488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1649977179
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_78
timestamp 1649977179
transform 1 0 8280 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_90
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_266
timestamp 1649977179
transform 1 0 25576 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1649977179
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_360
timestamp 1649977179
transform 1 0 34224 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_66
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_103
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_261
timestamp 1649977179
transform 1 0 25116 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_285
timestamp 1649977179
transform 1 0 27324 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_297
timestamp 1649977179
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1649977179
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_48
timestamp 1649977179
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_60
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_96
timestamp 1649977179
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1649977179
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_266
timestamp 1649977179
transform 1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_343
timestamp 1649977179
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_347
timestamp 1649977179
transform 1 0 33028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_358
timestamp 1649977179
transform 1 0 34040 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_261
timestamp 1649977179
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_284
timestamp 1649977179
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_296
timestamp 1649977179
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_10
timestamp 1649977179
transform 1 0 2024 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_22
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_38
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_199
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_211
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_265
timestamp 1649977179
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1649977179
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_55
timestamp 1649977179
transform 1 0 6164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_67
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1649977179
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_106
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_118
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1649977179
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_181
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_216
timestamp 1649977179
transform 1 0 20976 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_228
timestamp 1649977179
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_240
timestamp 1649977179
transform 1 0 23184 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_77
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_88
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_100
timestamp 1649977179
transform 1 0 10304 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_179
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_191
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_203
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_246
timestamp 1649977179
transform 1 0 23736 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_258
timestamp 1649977179
transform 1 0 24840 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1649977179
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1649977179
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_346
timestamp 1649977179
transform 1 0 32936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_358
timestamp 1649977179
transform 1 0 34040 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_285
timestamp 1649977179
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_291
timestamp 1649977179
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1649977179
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_14
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_308
timestamp 1649977179
transform 1 0 29440 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_320
timestamp 1649977179
transform 1 0 30544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_348
timestamp 1649977179
transform 1 0 33120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1649977179
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_11
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_17
timestamp 1649977179
transform 1 0 2668 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1649977179
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_106
timestamp 1649977179
transform 1 0 10856 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_118
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_130
timestamp 1649977179
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1649977179
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_286
timestamp 1649977179
transform 1 0 27416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_293
timestamp 1649977179
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_330
timestamp 1649977179
transform 1 0 31464 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_342
timestamp 1649977179
transform 1 0 32568 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1649977179
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1649977179
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_62
timestamp 1649977179
transform 1 0 6808 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_70
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_83
timestamp 1649977179
transform 1 0 8740 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1649977179
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_290
timestamp 1649977179
transform 1 0 27784 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_302
timestamp 1649977179
transform 1 0 28888 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_308
timestamp 1649977179
transform 1 0 29440 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_312
timestamp 1649977179
transform 1 0 29808 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_324
timestamp 1649977179
transform 1 0 30912 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_358
timestamp 1649977179
transform 1 0 34040 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_48
timestamp 1649977179
transform 1 0 5520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_120
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1649977179
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1649977179
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1649977179
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_329
timestamp 1649977179
transform 1 0 31372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_335
timestamp 1649977179
transform 1 0 31924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_342
timestamp 1649977179
transform 1 0 32568 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_351
timestamp 1649977179
transform 1 0 33396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1649977179
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_60
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_72
timestamp 1649977179
transform 1 0 7728 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_101
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_116
timestamp 1649977179
transform 1 0 11776 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_128
timestamp 1649977179
transform 1 0 12880 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_140
timestamp 1649977179
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_152
timestamp 1649977179
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1649977179
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1649977179
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1649977179
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_360
timestamp 1649977179
transform 1 0 34224 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_129
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1649977179
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_183
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_276
timestamp 1649977179
transform 1 0 26496 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_288
timestamp 1649977179
transform 1 0 27600 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_300
timestamp 1649977179
transform 1 0 28704 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_330
timestamp 1649977179
transform 1 0 31464 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_342
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_354
timestamp 1649977179
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1649977179
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_89
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_192
timestamp 1649977179
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_204
timestamp 1649977179
transform 1 0 19872 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1649977179
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_255
timestamp 1649977179
transform 1 0 24564 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1649977179
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1649977179
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1649977179
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_181
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1649977179
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_295
timestamp 1649977179
transform 1 0 28244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1649977179
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_312
timestamp 1649977179
transform 1 0 29808 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_324
timestamp 1649977179
transform 1 0 30912 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_336
timestamp 1649977179
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_348
timestamp 1649977179
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1649977179
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_321
timestamp 1649977179
transform 1 0 30636 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_325
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1649977179
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_360
timestamp 1649977179
transform 1 0 34224 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_207
timestamp 1649977179
transform 1 0 20148 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_219
timestamp 1649977179
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_231
timestamp 1649977179
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1649977179
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_315
timestamp 1649977179
transform 1 0 30084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_344
timestamp 1649977179
transform 1 0 32752 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_351
timestamp 1649977179
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_175
timestamp 1649977179
transform 1 0 17204 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1649977179
transform 1 0 17572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_189
timestamp 1649977179
transform 1 0 18492 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_195
timestamp 1649977179
transform 1 0 19044 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1649977179
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_212
timestamp 1649977179
transform 1 0 20608 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1649977179
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_360
timestamp 1649977179
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1649977179
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_207
timestamp 1649977179
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_219
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_231
timestamp 1649977179
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1649977179
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_315
timestamp 1649977179
transform 1 0 30084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_326
timestamp 1649977179
transform 1 0 31096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_334
timestamp 1649977179
transform 1 0 31832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_340
timestamp 1649977179
transform 1 0 32384 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1649977179
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 1649977179
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_92
timestamp 1649977179
transform 1 0 9568 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_98
timestamp 1649977179
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1649977179
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1649977179
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_325
timestamp 1649977179
transform 1 0 31004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_344
timestamp 1649977179
transform 1 0 32752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_356
timestamp 1649977179
transform 1 0 33856 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_71
timestamp 1649977179
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1649977179
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_88
timestamp 1649977179
transform 1 0 9200 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_117
timestamp 1649977179
transform 1 0 11868 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1649977179
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1649977179
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_326
timestamp 1649977179
transform 1 0 31096 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_351
timestamp 1649977179
transform 1 0 33396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_94
timestamp 1649977179
transform 1 0 9752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_101
timestamp 1649977179
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1649977179
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_301
timestamp 1649977179
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_307
timestamp 1649977179
transform 1 0 29348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1649977179
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_340
timestamp 1649977179
transform 1 0 32384 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_352
timestamp 1649977179
transform 1 0 33488 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_73
timestamp 1649977179
transform 1 0 7820 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_315
timestamp 1649977179
transform 1 0 30084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_327
timestamp 1649977179
transform 1 0 31188 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_349
timestamp 1649977179
transform 1 0 33212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp 1649977179
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_325
timestamp 1649977179
transform 1 0 31004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1649977179
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_267
timestamp 1649977179
transform 1 0 25668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_346
timestamp 1649977179
transform 1 0 32936 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1649977179
transform 1 0 33580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_360
timestamp 1649977179
transform 1 0 34224 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_257
timestamp 1649977179
transform 1 0 24748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_261
timestamp 1649977179
transform 1 0 25116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_286
timestamp 1649977179
transform 1 0 27416 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_293
timestamp 1649977179
transform 1 0 28060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1649977179
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1649977179
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 1649977179
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1649977179
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_303
timestamp 1649977179
transform 1 0 28980 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1649977179
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_360
timestamp 1649977179
transform 1 0 34224 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1649977179
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_117
timestamp 1649977179
transform 1 0 11868 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_122
timestamp 1649977179
transform 1 0 12328 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_134
timestamp 1649977179
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_147
timestamp 1649977179
transform 1 0 14628 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_159
timestamp 1649977179
transform 1 0 15732 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_171
timestamp 1649977179
transform 1 0 16836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_183
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_219
timestamp 1649977179
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_231
timestamp 1649977179
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1649977179
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 1649977179
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_283
timestamp 1649977179
transform 1 0 27140 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_290
timestamp 1649977179
transform 1 0 27784 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1649977179
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1649977179
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1649977179
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1649977179
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1649977179
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1649977179
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_286
timestamp 1649977179
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_298
timestamp 1649977179
transform 1 0 28520 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_310
timestamp 1649977179
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1649977179
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1649977179
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_345
timestamp 1649977179
transform 1 0 32844 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_356
timestamp 1649977179
transform 1 0 33856 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1649977179
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_105
timestamp 1649977179
transform 1 0 10764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_111
timestamp 1649977179
transform 1 0 11316 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_120
timestamp 1649977179
transform 1 0 12144 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1649977179
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_146
timestamp 1649977179
transform 1 0 14536 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_158
timestamp 1649977179
transform 1 0 15640 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_170
timestamp 1649977179
transform 1 0 16744 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_182
timestamp 1649977179
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1649977179
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_353
timestamp 1649977179
transform 1 0 33580 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1649977179
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_108
timestamp 1649977179
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_134
timestamp 1649977179
transform 1 0 13432 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_146
timestamp 1649977179
transform 1 0 14536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1649977179
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1649977179
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1649977179
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1649977179
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_269
timestamp 1649977179
transform 1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1649977179
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_302
timestamp 1649977179
transform 1 0 28888 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_314
timestamp 1649977179
transform 1 0 29992 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_326
timestamp 1649977179
transform 1 0 31096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1649977179
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_181
timestamp 1649977179
transform 1 0 17756 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_185
timestamp 1649977179
transform 1 0 18124 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1649977179
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_202
timestamp 1649977179
transform 1 0 19688 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_227
timestamp 1649977179
transform 1 0 21988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_239
timestamp 1649977179
transform 1 0 23092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_276
timestamp 1649977179
transform 1 0 26496 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_288
timestamp 1649977179
transform 1 0 27600 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 1649977179
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_329
timestamp 1649977179
transform 1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_334
timestamp 1649977179
transform 1 0 31832 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_346
timestamp 1649977179
transform 1 0 32936 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1649977179
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1649977179
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_207
timestamp 1649977179
transform 1 0 20148 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1649977179
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1649977179
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_358
timestamp 1649977179
transform 1 0 34040 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_185
timestamp 1649977179
transform 1 0 18124 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1649977179
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_285
timestamp 1649977179
transform 1 0 27324 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_290
timestamp 1649977179
transform 1 0 27784 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1649977179
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_330
timestamp 1649977179
transform 1 0 31464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1649977179
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_97
timestamp 1649977179
transform 1 0 10028 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_101
timestamp 1649977179
transform 1 0 10396 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 1649977179
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_287
timestamp 1649977179
transform 1 0 27508 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1649977179
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_321
timestamp 1649977179
transform 1 0 30636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1649977179
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_340
timestamp 1649977179
transform 1 0 32384 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_352
timestamp 1649977179
transform 1 0 33488 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1649977179
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_116
timestamp 1649977179
transform 1 0 11776 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_128
timestamp 1649977179
transform 1 0 12880 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_285
timestamp 1649977179
transform 1 0 27324 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_291
timestamp 1649977179
transform 1 0 27876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1649977179
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_99
timestamp 1649977179
transform 1 0 10212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_293
timestamp 1649977179
transform 1 0 28060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1649977179
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_177
timestamp 1649977179
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_199
timestamp 1649977179
transform 1 0 19412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_211
timestamp 1649977179
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_289
timestamp 1649977179
transform 1 0 27692 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_312
timestamp 1649977179
transform 1 0 29808 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_324
timestamp 1649977179
transform 1 0 30912 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_11
timestamp 1649977179
transform 1 0 2116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1649977179
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_181
timestamp 1649977179
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1649977179
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_294
timestamp 1649977179
transform 1 0 28152 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1649977179
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_65
timestamp 1649977179
transform 1 0 7084 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_70
timestamp 1649977179
transform 1 0 7544 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_82
timestamp 1649977179
transform 1 0 8648 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_94
timestamp 1649977179
transform 1 0 9752 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_106
timestamp 1649977179
transform 1 0 10856 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1649977179
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1649977179
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_184
timestamp 1649977179
transform 1 0 18032 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_209
timestamp 1649977179
transform 1 0 20332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1649977179
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_231
timestamp 1649977179
transform 1 0 22356 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_243
timestamp 1649977179
transform 1 0 23460 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_255
timestamp 1649977179
transform 1 0 24564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_267
timestamp 1649977179
transform 1 0 25668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_339
timestamp 1649977179
transform 1 0 32292 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_343
timestamp 1649977179
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_355
timestamp 1649977179
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_50
timestamp 1649977179
transform 1 0 5704 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_68
timestamp 1649977179
transform 1 0 7360 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_80
timestamp 1649977179
transform 1 0 8464 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_92
timestamp 1649977179
transform 1 0 9568 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_104
timestamp 1649977179
transform 1 0 10672 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_201
timestamp 1649977179
transform 1 0 19596 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_231
timestamp 1649977179
transform 1 0 22356 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_243
timestamp 1649977179
transform 1 0 23460 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_255
timestamp 1649977179
transform 1 0 24564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_267
timestamp 1649977179
transform 1 0 25668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_318
timestamp 1649977179
transform 1 0 30360 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_330
timestamp 1649977179
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_360
timestamp 1649977179
transform 1 0 34224 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_62
timestamp 1649977179
transform 1 0 6808 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1649977179
transform 1 0 18308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_220
timestamp 1649977179
transform 1 0 21344 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_228
timestamp 1649977179
transform 1 0 22080 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_297
timestamp 1649977179
transform 1 0 28428 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_341
timestamp 1649977179
transform 1 0 32476 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_347
timestamp 1649977179
transform 1 0 33028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_359
timestamp 1649977179
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1649977179
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1649977179
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_94
timestamp 1649977179
transform 1 0 9752 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_106
timestamp 1649977179
transform 1 0 10856 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1649977179
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1649977179
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_252
timestamp 1649977179
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_264
timestamp 1649977179
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1649977179
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_297
timestamp 1649977179
transform 1 0 28428 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_301
timestamp 1649977179
transform 1 0 28796 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_313
timestamp 1649977179
transform 1 0 29900 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_325
timestamp 1649977179
transform 1 0 31004 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 1649977179
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_57
timestamp 1649977179
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_69
timestamp 1649977179
transform 1 0 7452 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_76
timestamp 1649977179
transform 1 0 8096 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_113
timestamp 1649977179
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_125
timestamp 1649977179
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1649977179
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_164
timestamp 1649977179
transform 1 0 16192 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_169
timestamp 1649977179
transform 1 0 16652 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_176
timestamp 1649977179
transform 1 0 17296 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_183
timestamp 1649977179
transform 1 0 17940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_203
timestamp 1649977179
transform 1 0 19780 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_210
timestamp 1649977179
transform 1 0 20424 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_217
timestamp 1649977179
transform 1 0 21068 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_223
timestamp 1649977179
transform 1 0 21620 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_225
timestamp 1649977179
transform 1 0 21804 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_231
timestamp 1649977179
transform 1 0 22356 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_235
timestamp 1649977179
transform 1 0 22724 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1649977179
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_281
timestamp 1649977179
transform 1 0 26956 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_293
timestamp 1649977179
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1649977179
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_337
timestamp 1649977179
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_349
timestamp 1649977179
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1649977179
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 34868 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 34868 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 34868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 34868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 34868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 34868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 34868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 34868 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 34868 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _244_
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1649977179
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1649977179
transform 1 0 30544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1649977179
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1649977179
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _256_
timestamp 1649977179
transform 1 0 16928 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17204 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1649977179
transform 1 0 19504 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1649977179
transform 1 0 27508 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1649977179
transform 1 0 17020 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1649977179
transform -1 0 16192 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _263_
timestamp 1649977179
transform -1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1649977179
transform -1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1649977179
transform -1 0 5704 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1649977179
transform 1 0 24196 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1649977179
transform 1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1649977179
transform 1 0 22264 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _269_
timestamp 1649977179
transform -1 0 17756 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1649977179
transform 1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1649977179
transform 1 0 7820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1649977179
transform -1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1649977179
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _275_
timestamp 1649977179
transform 1 0 17940 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1649977179
transform 1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1649977179
transform 1 0 27140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1649977179
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1649977179
transform -1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1649977179
transform -1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _281_
timestamp 1649977179
transform -1 0 16928 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1649977179
transform -1 0 10488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1649977179
transform -1 0 28060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1649977179
transform -1 0 8464 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1649977179
transform 1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _288_
timestamp 1649977179
transform 1 0 19596 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1649977179
transform 1 0 28520 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1649977179
transform 1 0 29808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1649977179
transform 1 0 32384 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1649977179
transform -1 0 19964 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1649977179
transform 1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _294_
timestamp 1649977179
transform 1 0 17940 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1649977179
transform 1 0 25392 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1649977179
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1649977179
transform -1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1649977179
transform -1 0 3036 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _300_
timestamp 1649977179
transform -1 0 20148 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1649977179
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1649977179
transform 1 0 26128 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1649977179
transform -1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1649977179
transform 1 0 24840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _306_
timestamp 1649977179
transform 1 0 20056 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1649977179
transform -1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1649977179
transform -1 0 19964 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1649977179
transform -1 0 27784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _312_
timestamp 1649977179
transform 1 0 19136 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1649977179
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1649977179
transform 1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1649977179
transform 1 0 31556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1649977179
transform 1 0 32108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1649977179
transform -1 0 12328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1649977179
transform -1 0 16192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _319_
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1649977179
transform 1 0 31096 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1649977179
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1649977179
transform -1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1649977179
transform 1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _325_
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1649977179
transform -1 0 4968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1649977179
transform 1 0 17848 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1649977179
transform 1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _331_
timestamp 1649977179
transform -1 0 18768 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1649977179
transform 1 0 29072 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1649977179
transform -1 0 10396 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1649977179
transform -1 0 9292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1649977179
transform 1 0 22080 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1649977179
transform 1 0 27784 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _337_
timestamp 1649977179
transform -1 0 17572 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1649977179
transform 1 0 32476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1649977179
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1649977179
transform 1 0 32200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1649977179
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1649977179
transform 1 0 32476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _343_
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1649977179
transform -1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1649977179
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1649977179
transform 1 0 20148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1649977179
transform 1 0 27784 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _349_
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1649977179
transform -1 0 9200 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1649977179
transform 1 0 33120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1649977179
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1649977179
transform -1 0 32936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1649977179
transform -1 0 32936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _355_
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1649977179
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1649977179
transform 1 0 17480 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1649977179
transform -1 0 7544 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1649977179
transform -1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _361_
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1649977179
transform 1 0 33764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1649977179
transform -1 0 33580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1649977179
transform 1 0 33948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1649977179
transform -1 0 17664 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1649977179
transform 1 0 33120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _367_
timestamp 1649977179
transform -1 0 17572 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1649977179
transform -1 0 3128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1649977179
transform -1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1649977179
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484__2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _485__3
timestamp 1649977179
transform -1 0 18768 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _485_
timestamp 1649977179
transform 1 0 18400 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _486__4
timestamp 1649977179
transform 1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _486_
timestamp 1649977179
transform -1 0 8464 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _487__5
timestamp 1649977179
transform 1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _487_
timestamp 1649977179
transform 1 0 17480 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _488_
timestamp 1649977179
transform -1 0 7360 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _488__6
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489__7
timestamp 1649977179
transform -1 0 33120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _489_
timestamp 1649977179
transform 1 0 32292 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _490__8
timestamp 1649977179
transform -1 0 33212 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _490_
timestamp 1649977179
transform 1 0 32292 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _491_
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _491__9
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492__10
timestamp 1649977179
transform -1 0 33028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _492_
timestamp 1649977179
transform 1 0 32292 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _493__11
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _493_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _494__12
timestamp 1649977179
transform 1 0 28152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _494_
timestamp 1649977179
transform 1 0 29348 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _495__13
timestamp 1649977179
transform 1 0 19412 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _495_
timestamp 1649977179
transform 1 0 20056 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _496__14
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _496_
timestamp 1649977179
transform -1 0 13156 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _497__15
timestamp 1649977179
transform -1 0 29808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _497_
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _498__16
timestamp 1649977179
transform -1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _498_
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _499__17
timestamp 1649977179
transform -1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _499_
timestamp 1649977179
transform 1 0 32292 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _500__18
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _500_
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _501__19
timestamp 1649977179
transform -1 0 33120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _501_
timestamp 1649977179
transform 1 0 32292 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _502__20
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _502_
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _503__21
timestamp 1649977179
transform -1 0 33028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _503_
timestamp 1649977179
transform 1 0 32292 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _504__22
timestamp 1649977179
transform -1 0 28152 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _504_
timestamp 1649977179
transform 1 0 27876 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _505_
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _505__23
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _506__24
timestamp 1649977179
transform -1 0 22356 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _506_
timestamp 1649977179
transform 1 0 21988 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _507__25
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _507_
timestamp 1649977179
transform 1 0 8464 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _508__26
timestamp 1649977179
transform -1 0 10212 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _508_
timestamp 1649977179
transform 1 0 9844 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _509__27
timestamp 1649977179
transform -1 0 30084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _509_
timestamp 1649977179
transform 1 0 29716 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _510__28
timestamp 1649977179
transform -1 0 14536 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _510_
timestamp 1649977179
transform 1 0 14260 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _511__29
timestamp 1649977179
transform -1 0 18584 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _511_
timestamp 1649977179
transform 1 0 18216 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _512__30
timestamp 1649977179
transform -1 0 4508 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _512_
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _513__31
timestamp 1649977179
transform -1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _513_
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _514__32
timestamp 1649977179
transform 1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _514_
timestamp 1649977179
transform -1 0 8280 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _515__33
timestamp 1649977179
transform -1 0 31096 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _515_
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _516__34
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _516_
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _517__35
timestamp 1649977179
transform -1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _517_
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _518_
timestamp 1649977179
transform 1 0 30268 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _518__36
timestamp 1649977179
transform -1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_
timestamp 1649977179
transform 1 0 31464 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _519__37
timestamp 1649977179
transform 1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520__38
timestamp 1649977179
transform -1 0 12144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1649977179
transform 1 0 11776 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__39
timestamp 1649977179
transform -1 0 32752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1649977179
transform 1 0 32292 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _522__40
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _523__41
timestamp 1649977179
transform -1 0 32568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__42
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1649977179
transform 1 0 9108 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _525__43
timestamp 1649977179
transform -1 0 27416 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1649977179
transform 1 0 27048 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__44
timestamp 1649977179
transform -1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1649977179
transform 1 0 19320 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _527__45
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1649977179
transform 1 0 23920 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__46
timestamp 1649977179
transform -1 0 28612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1649977179
transform 1 0 28336 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _529__47
timestamp 1649977179
transform -1 0 20976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1649977179
transform 1 0 25208 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__48
timestamp 1649977179
transform -1 0 26404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531__49
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _532__50
timestamp 1649977179
transform 1 0 26220 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _533__51
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _534__52
timestamp 1649977179
transform -1 0 27508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1649977179
transform 1 0 27232 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _535__53
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _536__54
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__55
timestamp 1649977179
transform -1 0 3128 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1649977179
transform 1 0 2760 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1649977179
transform 1 0 27784 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _538__56
timestamp 1649977179
transform -1 0 28152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539__57
timestamp 1649977179
transform -1 0 25760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _540__58
timestamp 1649977179
transform -1 0 32384 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1649977179
transform 1 0 31832 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__59
timestamp 1649977179
transform 1 0 20148 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1649977179
transform -1 0 21160 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__60
timestamp 1649977179
transform -1 0 33028 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1649977179
transform 1 0 32292 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _543__61
timestamp 1649977179
transform -1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1649977179
transform 1 0 29716 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__62
timestamp 1649977179
transform -1 0 30084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _545__63
timestamp 1649977179
transform -1 0 28796 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1649977179
transform 1 0 28428 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1649977179
transform 1 0 19412 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__64
timestamp 1649977179
transform -1 0 19780 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _547__65
timestamp 1649977179
transform -1 0 29992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__66
timestamp 1649977179
transform -1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1649977179
transform 1 0 7636 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _549__67
timestamp 1649977179
transform -1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1649977179
transform 1 0 27508 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__68
timestamp 1649977179
transform -1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1649977179
transform 1 0 9936 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _551__69
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _551_
timestamp 1649977179
transform -1 0 8096 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _552_
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _552__70
timestamp 1649977179
transform -1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _553__71
timestamp 1649977179
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _553_
timestamp 1649977179
transform -1 0 7176 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _554_
timestamp 1649977179
transform 1 0 27140 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _554__72
timestamp 1649977179
transform -1 0 27784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _555_
timestamp 1649977179
transform 1 0 25300 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _555__73
timestamp 1649977179
transform -1 0 25576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _556__74
timestamp 1649977179
transform -1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _556_
timestamp 1649977179
transform 1 0 25392 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _557__75
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _557_
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _558__76
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _558_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _559__77
timestamp 1649977179
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _559_
timestamp 1649977179
transform 1 0 27508 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _560__78
timestamp 1649977179
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _560_
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _561__79
timestamp 1649977179
transform -1 0 22724 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _561_
timestamp 1649977179
transform 1 0 22356 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _562__80
timestamp 1649977179
transform -1 0 8096 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _562_
timestamp 1649977179
transform 1 0 7820 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _563__81
timestamp 1649977179
transform -1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _563_
timestamp 1649977179
transform 1 0 24564 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _564__82
timestamp 1649977179
transform -1 0 5244 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _564_
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _565__83
timestamp 1649977179
transform -1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _565_
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _566__84
timestamp 1649977179
transform 1 0 15916 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _566_
timestamp 1649977179
transform 1 0 16376 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _567__85
timestamp 1649977179
transform -1 0 17940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _567_
timestamp 1649977179
transform 1 0 16928 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _568__86
timestamp 1649977179
transform -1 0 29808 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _568_
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _569__87
timestamp 1649977179
transform -1 0 27876 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _569_
timestamp 1649977179
transform 1 0 27600 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _570__88
timestamp 1649977179
transform 1 0 20792 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _570_
timestamp 1649977179
transform -1 0 21344 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _571_
timestamp 1649977179
transform 1 0 30912 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _571__89
timestamp 1649977179
transform -1 0 31648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _572__90
timestamp 1649977179
transform -1 0 31556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _572_
timestamp 1649977179
transform 1 0 31280 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _573__91
timestamp 1649977179
transform 1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _573_
timestamp 1649977179
transform -1 0 9752 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _574__92
timestamp 1649977179
transform -1 0 31464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _574_
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _575__93
timestamp 1649977179
transform -1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _575_
timestamp 1649977179
transform 1 0 10212 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _576__94
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _576_
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _577__95
timestamp 1649977179
transform -1 0 5520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _577_
timestamp 1649977179
transform 1 0 5152 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _578__96
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _578_
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _579__97
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _579_
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _580_
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _580__98
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _581__99
timestamp 1649977179
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _581_
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _582__100
timestamp 1649977179
transform -1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _582_
timestamp 1649977179
transform 1 0 2760 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _583_
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _583__101
timestamp 1649977179
transform -1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _584__102
timestamp 1649977179
transform -1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _584_
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _585__103
timestamp 1649977179
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _585_
timestamp 1649977179
transform 1 0 17572 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _586__104
timestamp 1649977179
transform -1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _586_
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _587_
timestamp 1649977179
transform -1 0 34224 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _587__105
timestamp 1649977179
transform 1 0 33764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _588__106
timestamp 1649977179
transform 1 0 16744 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _588_
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _589__107
timestamp 1649977179
transform 1 0 33764 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _589_
timestamp 1649977179
transform -1 0 34224 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _590__108
timestamp 1649977179
transform 1 0 33580 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _590_
timestamp 1649977179
transform -1 0 34224 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _591__109
timestamp 1649977179
transform 1 0 33764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _591_
timestamp 1649977179
transform -1 0 34224 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 35904
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 35988 800 36228 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 11582 0 11694 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 18666 41200 18778 42000 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal3 s 0 38708 800 38948 0 FreeSans 960 0 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 35200 35988 36000 36228 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18022 0 18134 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 11582 41200 11694 42000 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 35200 37348 36000 37588 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 35200 6068 36000 6308 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 5142 41200 5254 42000 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 6430 41200 6542 42000 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 33478 0 33590 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 0 12188 800 12428 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 0 22388 800 22628 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 0 14908 800 15148 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 35200 15588 36000 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 4498 41200 4610 42000 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 1922 41200 2034 42000 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 28970 0 29082 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 28326 0 28438 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 35200 11508 36000 11748 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 35410 41200 35522 42000 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 12870 0 12982 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 35200 18308 36000 18548 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 0 34628 800 34868 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 23818 0 23930 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 0 20348 800 20588 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 26394 41200 26506 42000 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 30902 41200 31014 42000 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 35200 27148 36000 27388 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 31546 41200 31658 42000 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 19310 41200 19422 42000 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 35200 26468 36000 26708 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 35200 40068 36000 40308 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 0 23748 800 23988 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 0 16268 800 16508 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 35200 29188 36000 29428 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 3210 41200 3322 42000 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal3 s 0 13548 800 13788 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal3 s 35200 25108 36000 25348 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal3 s 35200 14228 36000 14468 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal3 s 35200 13548 36000 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 7718 41200 7830 42000 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal3 s 35200 4708 36000 4948 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 10294 0 10406 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 25106 41200 25218 42000 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 8362 41200 8474 42000 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 30258 0 30370 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal3 s 35200 19668 36000 19908 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal3 s 0 40748 800 40988 0 FreeSans 960 0 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 3854 0 3966 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 16090 41200 16202 42000 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 17378 41200 17490 42000 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal3 s 35200 628 36000 868 0 FreeSans 960 0 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal3 s 35200 33268 36000 33508 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 19954 41200 20066 42000 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 32834 0 32946 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal3 s 35200 27828 36000 28068 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 28970 41200 29082 42000 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal3 s 0 41428 800 41668 0 FreeSans 960 0 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal3 s 0 18988 800 19228 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal3 s 35200 1988 36000 2228 0 FreeSans 960 0 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 5786 41200 5898 42000 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal3 s 0 8788 800 9028 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal3 s 0 14228 800 14468 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 19954 0 20066 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal3 s 35200 3348 36000 3588 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal3 s 0 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal3 s 35200 16948 36000 17188 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 7074 41200 7186 42000 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 8362 0 8474 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal3 s 35200 39388 36000 39628 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal3 s 35200 24428 36000 24668 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal3 s 0 1988 800 2228 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal3 s 0 5388 800 5628 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 30902 0 31014 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal3 s 35200 33948 36000 34188 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal3 s 0 31908 800 32148 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal3 s 35200 23748 36000 23988 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 32834 41200 32946 42000 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal3 s 35200 -52 36000 188 0 FreeSans 960 0 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 22530 41200 22642 42000 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 28326 41200 28438 42000 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal3 s 0 31228 800 31468 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 24462 0 24574 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal3 s 35200 20348 36000 20588 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 21242 0 21354 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 25750 41200 25862 42000 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal3 s 0 4028 800 4268 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 27038 41200 27150 42000 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 13514 0 13626 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal3 s 35200 4028 36000 4268 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 5142 0 5254 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal3 s 0 10828 800 11068 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal3 s 0 36668 800 36908 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal3 s 35200 8788 36000 9028 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal3 s 35200 34628 36000 34868 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal3 s 35200 32588 36000 32828 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 9006 41200 9118 42000 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal3 s 35200 38028 36000 38268 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal3 s 0 33948 800 34188 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal3 s 35200 25788 36000 26028 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 14802 41200 14914 42000 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 34122 41200 34234 42000 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal3 s 0 15588 800 15828 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 14802 0 14914 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal3 s 35200 9468 36000 9708 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 16734 0 16846 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 35200 7428 36000 7668 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 0 29188 800 29428 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 26394 0 26506 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 9650 41200 9762 42000 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 21242 41200 21354 42000 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 15446 41200 15558 42000 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 34122 0 34234 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 10938 41200 11050 42000 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 15446 0 15558 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 0 28508 800 28748 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 34766 41200 34878 42000 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 35200 10148 36000 10388 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 0 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 0 29868 800 30108 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 35200 5388 36000 5628 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 0 25788 800 26028 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal3 s 0 39388 800 39628 0 FreeSans 960 0 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 9006 0 9118 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 0 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 29614 0 29726 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 0 24428 800 24668 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 30258 41200 30370 42000 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 35200 22388 36000 22628 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 12226 41200 12338 42000 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 0 17628 800 17868 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 12870 41200 12982 42000 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 0 27148 800 27388 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal tristate
flabel metal3 s 35200 12188 36000 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal tristate
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal tristate
flabel metal3 s 35200 38708 36000 38948 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal tristate
flabel metal2 s 634 41200 746 42000 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal tristate
flabel metal2 s 18022 41200 18134 42000 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal tristate
flabel metal3 s 0 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal tristate
flabel metal3 s 35200 16268 36000 16508 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal tristate
flabel metal3 s 35200 31228 36000 31468 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal tristate
flabel metal2 s 1278 41200 1390 42000 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal tristate
flabel metal3 s 35200 23068 36000 23308 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal tristate
flabel metal3 s 0 35308 800 35548 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal tristate
flabel metal3 s 0 8108 800 8348 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal tristate
flabel metal3 s 35200 36668 36000 36908 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal tristate
flabel metal2 s 20598 41200 20710 42000 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal tristate
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal tristate
flabel metal3 s 35200 17628 36000 17868 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal tristate
flabel metal3 s 0 2668 800 2908 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal tristate
flabel metal3 s 35200 6748 36000 6988 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal tristate
flabel metal3 s 0 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal tristate
flabel metal2 s 34766 0 34878 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal tristate
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal tristate
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal tristate
flabel metal3 s 35200 12868 36000 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal tristate
flabel metal3 s 35200 40748 36000 40988 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal tristate
flabel metal3 s 0 7428 800 7668 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal tristate
flabel metal2 s 35410 0 35522 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal tristate
flabel metal2 s 2566 0 2678 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal tristate
flabel metal3 s 35200 18988 36000 19228 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal tristate
flabel metal2 s 634 0 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal tristate
flabel metal3 s 35200 31908 36000 32148 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal tristate
flabel metal2 s 33478 41200 33590 42000 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal tristate
flabel metal3 s 35200 2668 36000 2908 0 FreeSans 960 0 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 32190 41200 32302 42000 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 0 21708 800 21948 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 0 23068 800 23308 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 23174 0 23286 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 27682 0 27794 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 0 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s -10 41200 102 42000 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 14158 41200 14270 42000 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 0 21028 800 21268 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 7074 0 7186 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 1922 0 2034 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 21886 41200 21998 42000 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 13514 41200 13626 42000 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 19310 0 19422 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 27682 41200 27794 42000 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 35200 10828 36000 11068 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 0 30548 800 30788 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 35200 30548 36000 30788 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 7718 0 7830 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 14158 0 14270 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 35200 29868 36000 30108 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 21886 0 21998 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 24462 41200 24574 42000 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 23818 41200 23930 42000 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 0 38028 800 38268 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 2566 41200 2678 42000 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 0 9468 800 9708 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 0 32588 800 32828 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 5168 2128 5488 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 13616 2128 13936 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 22064 2128 22384 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 30512 2128 30832 39760 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 9392 2128 9712 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 17840 2128 18160 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal4 s 26288 2128 26608 39760 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 35200 21028 36000 21268 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36000 42000
<< end >>
